library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity top is
port (
    clkin_50                    : in    std_logic--;
);
end entity;

architecture arch of top is

begin

end architecture;

library ieee;
use ieee.std_logic_1164.all;

-- 8b10b decoder
-- https://en.wikipedia.org/wiki/8b/10b_encoding
entity dec_8b10b is
    port (
        -- input 10-bit data (8b10b encoded)
        datain  :   in  std_logic_vector(9 downto 0);
        -- input disparity
        dispin  :   in  std_logic;
        -- output data (K bit & 8 data bits)
        dataout :   out std_logic_vector(8 downto 0);
        -- output disparity
        dispout :   out std_logic;
        -- disparity error
        disperr :   out std_logic;
        -- error if invalid code
        err     :   out std_logic--;
    );
end entity;

architecture arch of dec_8b10b is

    -- control (K) symbol
    signal K : std_logic;

    -- 6-bit group --
    -- disp & 6 bits in
    signal g6sel : std_logic_vector(6 downto 0);
    -- err & disperr & disp & 5 bits out
    signal g6 : std_logic_vector(7 downto 0);

    signal K28, Kx7 : std_logic;

    -- 4-bit group --
    -- K.28 & disp & 4 bits in
    signal g4sel : std_logic_vector(5 downto 0);
    -- err & disperr & disp & 3 bits out
    signal g4 : std_logic_vector(5 downto 0);

begin

    K28 <= work.util.to_std_logic( datain(5 downto 0) = "111100" or datain(5 downto 0) = "000011" );
    Kx7 <= work.util.to_std_logic( ( datain(9 downto 6) = "0001" or datain(9 downto 6) = "1110" ) and (
        g6(4 downto 0) = "10111" or -- D.23
        g6(4 downto 0) = "11011" or -- D.27
        g6(4 downto 0) = "11101" or -- D.29
        g6(4 downto 0) = "11110" ) -- D.30
    );
    K <= '0';

    -- disp & 6 bits in
    g6sel <= dispin & datain(5 downto 0);
    -- err & disperr & disp & 5 bits out
    with g6sel select g6 <=
        '0' & '0' & '1' & "00000" when '0' & "111001",
        '0' & '0' & '0' & "00000" when '1' & "000110",
        '0' & '0' & '1' & "00001" when '0' & "101110",
        '0' & '0' & '0' & "00001" when '1' & "010001",
        '0' & '0' & '1' & "00010" when '0' & "101101",
        '0' & '0' & '0' & "00010" when '1' & "010010",
        '0' & '0' & '0' & "00011" when '0' & "100011",
        '0' & '0' & '1' & "00011" when '1' & "100011",
        '0' & '0' & '1' & "00100" when '0' & "101011",
        '0' & '0' & '0' & "00100" when '1' & "010100",
        '0' & '0' & '0' & "00101" when '0' & "100101",
        '0' & '0' & '1' & "00101" when '1' & "100101",
        '0' & '0' & '0' & "00110" when '0' & "100110",
        '0' & '0' & '1' & "00110" when '1' & "100110",
        '0' & '0' & '0' & "00111" when '0' & "000111", -- D.07
        '0' & '0' & '1' & "00111" when '1' & "111000", -- D.07
        '0' & '0' & '1' & "01000" when '0' & "100111",
        '0' & '0' & '0' & "01000" when '1' & "011000",
        '0' & '0' & '0' & "01001" when '0' & "101001",
        '0' & '0' & '1' & "01001" when '1' & "101001",
        '0' & '0' & '0' & "01010" when '0' & "101010",
        '0' & '0' & '1' & "01010" when '1' & "101010",
        '0' & '0' & '0' & "01011" when '0' & "001011",
        '0' & '0' & '1' & "01011" when '1' & "001011", -- D.11.A7
        '0' & '0' & '0' & "01100" when '0' & "101100",
        '0' & '0' & '1' & "01100" when '1' & "101100",
        '0' & '0' & '0' & "01101" when '0' & "001101",
        '0' & '0' & '1' & "01101" when '1' & "001101", -- D.13.A7
        '0' & '0' & '0' & "01110" when '0' & "001110",
        '0' & '0' & '1' & "01110" when '1' & "001110", -- D.14.A7
        '0' & '0' & '1' & "01111" when '0' & "111010",
        '0' & '0' & '0' & "01111" when '1' & "000101",
        '0' & '0' & '1' & "10000" when '0' & "110110",
        '0' & '0' & '0' & "10000" when '1' & "001001",
        '0' & '0' & '0' & "10001" when '0' & "110001", -- D.17.A7
        '0' & '0' & '1' & "10001" when '1' & "110001",
        '0' & '0' & '0' & "10010" when '0' & "110010", -- D.18.A7
        '0' & '0' & '1' & "10010" when '1' & "110010",
        '0' & '0' & '0' & "10011" when '0' & "010011",
        '0' & '0' & '1' & "10011" when '1' & "010011",
        '0' & '0' & '0' & "10100" when '0' & "110100", -- D.20.A7
        '0' & '0' & '1' & "10100" when '1' & "110100",
        '0' & '0' & '0' & "10101" when '0' & "010101",
        '0' & '0' & '1' & "10101" when '1' & "010101",
        '0' & '0' & '0' & "10110" when '0' & "010110",
        '0' & '0' & '1' & "10110" when '1' & "010110",
        '0' & '0' & '1' & "10111" when '0' & "010111",
        '0' & '0' & '0' & "10111" when '1' & "101000",
        '0' & '0' & '1' & "11000" when '0' & "110011",
        '0' & '0' & '0' & "11000" when '1' & "001100",
        '0' & '0' & '0' & "11001" when '0' & "011001",
        '0' & '0' & '1' & "11001" when '1' & "011001",
        '0' & '0' & '0' & "11010" when '0' & "011010",
        '0' & '0' & '1' & "11010" when '1' & "011010",
        '0' & '0' & '1' & "11011" when '0' & "011011",
        '0' & '0' & '0' & "11011" when '1' & "100100",
        '0' & '0' & '0' & "11100" when '0' & "011100", -- D.28
        '0' & '0' & '1' & "11100" when '1' & "011100", -- D.28
        '0' & '0' & '1' & "11100" when '0' & "111100", -- K.28
        '0' & '0' & '0' & "11100" when '1' & "000011", -- K.28
        '0' & '0' & '1' & "11101" when '0' & "011101",
        '0' & '0' & '0' & "11101" when '1' & "100010",
        '0' & '0' & '1' & "11110" when '0' & "011110",
        '0' & '0' & '0' & "11110" when '1' & "100001",
        '0' & '0' & '1' & "11111" when '0' & "110101",
        '0' & '0' & '0' & "11111" when '1' & "001010",
        -- invalid disparity
        '0' & '1' & '1' & "00000" when '1' & "111001",
        '0' & '1' & '0' & "00000" when '0' & "000110",
        '0' & '1' & '1' & "00001" when '1' & "101110",
        '0' & '1' & '0' & "00001" when '0' & "010001",
        '0' & '1' & '1' & "00010" when '1' & "101101",
        '0' & '1' & '0' & "00010" when '0' & "010010",
        '0' & '1' & '1' & "00100" when '1' & "101011",
        '0' & '1' & '0' & "00100" when '0' & "010100",
        '0' & '1' & '1' & "01000" when '1' & "100111",
        '0' & '1' & '0' & "01000" when '0' & "011000",
        '0' & '1' & '1' & "01111" when '1' & "111010",
        '0' & '1' & '0' & "01111" when '0' & "000101",
        '0' & '1' & '1' & "10000" when '1' & "110110",
        '0' & '1' & '0' & "10000" when '0' & "001001",
        '0' & '1' & '1' & "10111" when '1' & "010111",
        '0' & '1' & '0' & "10111" when '0' & "101000",
        '0' & '1' & '1' & "11000" when '1' & "110011",
        '0' & '1' & '0' & "11000" when '0' & "001100",
        '0' & '1' & '1' & "11011" when '1' & "011011",
        '0' & '1' & '0' & "11011" when '0' & "100100",
        '0' & '1' & '1' & "11100" when '1' & "111100", -- K.28
        '0' & '1' & '0' & "11100" when '0' & "000011", -- K.28
        '0' & '1' & '1' & "11101" when '1' & "011101",
        '0' & '1' & '0' & "11101" when '0' & "100010",
        '0' & '1' & '1' & "11110" when '1' & "011110",
        '0' & '1' & '0' & "11110" when '0' & "100001",
        '0' & '1' & '1' & "11111" when '1' & "110101",
        '0' & '1' & '0' & "11111" when '0' & "001010",
        --
        '0' & '1' & '1' & "00111" when '1' & "000111", -- D.07
        '0' & '1' & '0' & "00111" when '0' & "111000", -- D.07
        -- invalid code
        '1' & '0' & '1' & "XXXXX" when '0' & "001111",
        '1' & '0' & '0' & "XXXXX" when '1' & "110000",
        -- invalid code and disparity
        '1' & '1' & '1' & "XXXXX" when '1' & "001111",
        '1' & '1' & '0' & "XXXXX" when '0' & "110000",
        '1' & '1' & '1' & "XXXXX" when '0' & "111111",
        '1' & '1' & '0' & "XXXXX" when '1' & "000000",
        '1' & '1' & '1' & "XXXXX" when '1' & "111111",
        '1' & '1' & '0' & "XXXXX" when '0' & "000000",
        '1' & '1' & '1' & "XXXXX" when '0' & "111110",
        '1' & '1' & '0' & "XXXXX" when '1' & "000001",
        '1' & '1' & '1' & "XXXXX" when '1' & "111110",
        '1' & '1' & '0' & "XXXXX" when '0' & "000001",
        '1' & '1' & '1' & "XXXXX" when '0' & "111101",
        '1' & '1' & '0' & "XXXXX" when '1' & "000010",
        '1' & '1' & '1' & "XXXXX" when '1' & "111101",
        '1' & '1' & '0' & "XXXXX" when '0' & "000010",
        '1' & '1' & '1' & "XXXXX" when '0' & "111011",
        '1' & '1' & '0' & "XXXXX" when '1' & "000100",
        '1' & '1' & '1' & "XXXXX" when '1' & "111011",
        '1' & '1' & '0' & "XXXXX" when '0' & "000100",
        '1' & '1' & '1' & "XXXXX" when '0' & "110111",
        '1' & '1' & '0' & "XXXXX" when '1' & "001000",
        '1' & '1' & '1' & "XXXXX" when '1' & "110111",
        '1' & '1' & '0' & "XXXXX" when '0' & "001000",
        '1' & '1' & '1' & "XXXXX" when '0' & "101111",
        '1' & '1' & '0' & "XXXXX" when '1' & "010000",
        '1' & '1' & '1' & "XXXXX" when '1' & "101111",
        '1' & '1' & '0' & "XXXXX" when '0' & "010000",
        '1' & '1' & '1' & "XXXXX" when '0' & "011111",
        '1' & '1' & '0' & "XXXXX" when '1' & "100000",
        '1' & '1' & '1' & "XXXXX" when '1' & "011111",
        '1' & '1' & '0' & "XXXXX" when '0' & "100000",
        '1' & '1' & '0' & "XXXXX" when others;

    -- K.28 & disp & 4 bits in
    g4sel <= K28 & g6(5) & datain(9 downto 6);
    -- err & disperr & disp & 3 bits out
    with g4sel select g4 <=
        '0' & '0' & '1' & "000" when '0' & '0' & "1101", -- D.x.0
        '0' & '0' & '0' & "000" when '0' & '1' & "0010", -- D.x.0
        '0' & '0' & '0' & "001" when '0' & '0' & "1001", -- D.x.1
        '0' & '0' & '1' & "001" when '0' & '1' & "1001", -- D.x.1
        '0' & '0' & '0' & "010" when '0' & '0' & "1010", -- D.x.2
        '0' & '0' & '1' & "010" when '0' & '1' & "1010", -- D.x.2
        '0' & '0' & '0' & "011" when '0' & '0' & "0011", -- D.x.3
        '0' & '0' & '1' & "011" when '0' & '1' & "1100", -- D.x.3
        '0' & '0' & '1' & "100" when '0' & '0' & "1011", -- D.x.4
        '0' & '0' & '0' & "100" when '0' & '1' & "0100", -- D.x.4
        '0' & '0' & '0' & "101" when '0' & '0' & "0101", -- D.x.5
        '0' & '0' & '1' & "101" when '0' & '1' & "0101", -- D.x.5
        '0' & '0' & '0' & "110" when '0' & '0' & "0110", -- D.x.6
        '0' & '0' & '1' & "110" when '0' & '1' & "0110", -- D.x.6
        '0' & '0' & '1' & "111" when '0' & '0' & "0111", -- D.x.P7
        '0' & '0' & '0' & "111" when '0' & '1' & "1000", -- D.x.P7
        '0' & '0' & '1' & "111" when '0' & '0' & "1110", -- D.x.A7, K.x.7
        '0' & '0' & '0' & "111" when '0' & '1' & "0001", -- D.x.A7, K.x.7
        '0' & '0' & '1' & "000" when '1' & '0' & "1101", -- K.28.0
        '0' & '0' & '0' & "000" when '1' & '1' & "0010", -- K.28.0
        '0' & '0' & '0' & "001" when '1' & '0' & "0110", -- K.28.1
        '0' & '0' & '1' & "001" when '1' & '1' & "1001", -- K.28.1
        '0' & '0' & '0' & "010" when '1' & '0' & "0101", -- K.28.2
        '0' & '0' & '1' & "010" when '1' & '1' & "1010", -- K.28.2
        '0' & '0' & '0' & "011" when '1' & '0' & "0011", -- K.28.3
        '0' & '0' & '1' & "011" when '1' & '1' & "1100", -- K.28.3
        '0' & '0' & '1' & "100" when '1' & '0' & "1011", -- K.28.4
        '0' & '0' & '0' & "100" when '1' & '1' & "0100", -- K.28.4
        '0' & '0' & '0' & "101" when '1' & '0' & "1010", -- K.28.5
        '0' & '0' & '1' & "101" when '1' & '1' & "0101", -- K.28.5
        '0' & '0' & '0' & "110" when '1' & '0' & "1001", -- K.28.6
        '0' & '0' & '1' & "110" when '1' & '1' & "0110", -- K.28.6
        '0' & '0' & '1' & "111" when '1' & '0' & "1110", -- K.28.7
        '0' & '0' & '0' & "111" when '1' & '1' & "0001", -- K.28.7
        -- invalid disparity
        '0' & '1' & '1' & "000" when '0' & '1' & "1101", -- D.x.0
        '0' & '1' & '0' & "000" when '0' & '0' & "0010", -- D.x.0
        '0' & '1' & '1' & "000" when '1' & '1' & "1101", -- K.28.0
        '0' & '1' & '0' & "000" when '1' & '0' & "0010", -- K.28.0
        '0' & '1' & '1' & "100" when '0' & '1' & "1011", -- D.x.4
        '0' & '1' & '0' & "100" when '0' & '0' & "0100", -- D.x.4
        '0' & '1' & '1' & "100" when '1' & '1' & "1011", -- K.28.4
        '0' & '1' & '0' & "100" when '1' & '0' & "0100", -- K.28.4
        '0' & '1' & '1' & "111" when '0' & '1' & "0111", -- D.x.P7
        '0' & '1' & '0' & "111" when '0' & '0' & "1000", -- D.x.P7
        '0' & '1' & '1' & "111" when '0' & '1' & "1110", -- D.x.A7
        '0' & '1' & '0' & "111" when '0' & '0' & "0001", -- D.x.A7
        '0' & '1' & '1' & "111" when '1' & '1' & "1110", -- K.28.7
        '0' & '1' & '0' & "111" when '1' & '0' & "0001", -- K.28.7
        --
        '0' & '1' & '1' & "011" when '0' & '1' & "0011", -- D.x.3
        '0' & '1' & '0' & "011" when '0' & '0' & "1100", -- D.x.3
        '0' & '1' & '1' & "011" when '1' & '1' & "0011", -- K.28.3
        '0' & '1' & '0' & "011" when '1' & '0' & "1100", -- K.28.3
        -- invalid code
        '1' & '0' & '1' & "111" when '1' & '0' & "0111", -- D.x.P7
        '1' & '0' & '0' & "111" when '1' & '1' & "1000", -- D.x.P7
        '1' & '1' & '1' & "111" when '1' & '1' & "0111", -- D.x.P7
        '1' & '1' & '0' & "111" when '1' & '0' & "1000", -- D.x.P7
        -- invalid code and disparity
        '1' & '1' & '1' & "XXX" when '0' & '0' & "1111",
        '1' & '1' & '0' & "XXX" when '0' & '1' & "0000",
        '1' & '1' & '1' & "XXX" when '0' & '1' & "1111",
        '1' & '1' & '0' & "XXX" when '0' & '0' & "0000",
        '1' & '1' & '1' & "XXX" when '1' & '0' & "1111",
        '1' & '1' & '0' & "XXX" when '1' & '1' & "0000",
        '1' & '1' & '1' & "XXX" when '1' & '1' & "1111",
        '1' & '1' & '0' & "XXX" when '1' & '0' & "0000",
        '1' & '1' & '0' & "XXX" when others;

    dataout(4 downto 0) <= g6(4 downto 0);
    dataout(7 downto 5) <= g4(2 downto 0);
    dataout(8) <= K28 or Kx7;
    dispout <= g4(3);

    disperr <= g6(6) or g4(4);

    err <=
       work.util.to_std_logic(
           ( g6(4 downto 0) = "10001" or g6(4 downto 0) = "10010" or g6(4 downto 0) = "10100" )
           and g4(2 downto 0) = "111"
           and datain(9 downto 6) /= "1110" -- D.x.A7
       ) or
       work.util.to_std_logic(
           ( g6(4 downto 0) = "01110" or g6(4 downto 0) = "01101" or g6(4 downto 0) = "01011" )
           and g4(2 downto 0) = "111"
           and datain(9 downto 6) /= "0001" -- D.x.A7
       ) or
       g6(7) or g4(5);

end architecture;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package altera is

end package;

package body altera is

end package body;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tb_8b10b is
end entity;

architecture arch of tb_8b10b is

    type data_enc_t is array (natural range <>) of std_logic_vector(0 to 21);
    signal data_enc : data_enc_t(0 to 1023) := (
        -- dispin, k, d8, dispout, d10, err
        "0000000000000101110010","1000000000111010001100","0000000001000101011100","1000000001111010100010","0000000010000101011010","1000000010111010100100","0000000011111011000110","1000000011000101000110","0000000100000101010110","1000000100111010101000","0000000101111011001010","1000000101000101001010","0000000110111011001100","1000000110000101001100","0000000111111010001110","1000000111000101110000","0000001000000101001110","1000001000111010110000","0000001001111011010010","1000001001000101010010","0000001010111011010100","1000001010000101010100","0000001011111010010110","1000001011000100010110","0000001100111011011000","1000001100000101011000","0000001101111010011010","1000001101000100011010","0000001110111010011100","1000001110000100011100","0000001111000101110100","1000001111111010001010","0000010000000101101100","1000010000111010010010","0000010001111011100010","1000010001000101100010","0000010010111011100100","1000010010000101100100","0000010011111010100110","1000010011000100100110","0000010100111011101000","1000010100000101101000","0000010101111010101010","1000010101000100101010","0000010110111010101100","1000010110000100101100","0000010111000100101110","1000010111111011010000","0000011000000101100110","1000011000111010011000","0000011001111010110010","1000011001000100110010","0000011010111010110100","1000011010000100110100","0000011011000100110110","1000011011111011001000","0000011100111010111000","1000011100000100111000","0000011101000100111010","1000011101111011000100","0000011110000100111100","1000011110111011000010","0000011111000101101010","1000011111111010010100","0000100000110011110010","1000100000010010001100","0000100001110011011100","1000100001010010100010","0000100010110011011010","1000100010010010100100","0000100011010011000110","1000100011110011000110","0000100100110011010110","1000100100010010101000","0000100101010011001010","1000100101110011001010","0000100110010011001100","1000100110110011001100","0000100111010010001110","1000100111110011110000","0000101000110011001110","1000101000010010110000","0000101001010011010010","1000101001110011010010","0000101010010011010100","1000101010110011010100","0000101011010010010110","1000101011110010010110","0000101100010011011000","1000101100110011011000","0000101101010010011010","1000101101110010011010","0000101110010010011100","1000101110110010011100","0000101111110011110100","1000101111010010001010","0000110000110011101100","1000110000010010010010","0000110001010011100010","1000110001110011100010","0000110010010011100100","1000110010110011100100","0000110011010010100110","1000110011110010100110","0000110100010011101000","1000110100110011101000","0000110101010010101010","1000110101110010101010","0000110110010010101100","1000110110110010101100","0000110111110010101110","1000110111010011010000","0000111000110011100110","1000111000010010011000","0000111001010010110010","1000111001110010110010","0000111010010010110100","1000111010110010110100","0000111011110010110110","1000111011010011001000","0000111100010010111000","1000111100110010111000","0000111101110010111010","1000111101010011000100","0000111110110010111100","1000111110010011000010","0000111111110011101010","1000111111010010010100","0001000000110101110010","1001000000010100001100","0001000001110101011100","1001000001010100100010","0001000010110101011010","1001000010010100100100","0001000011010101000110","1001000011110101000110","0001000100110101010110","1001000100010100101000","0001000101010101001010","1001000101110101001010","0001000110010101001100","1001000110110101001100","0001000111010100001110","1001000111110101110000","0001001000110101001110","1001001000010100110000","0001001001010101010010","1001001001110101010010","0001001010010101010100","1001001010110101010100","0001001011010100010110","1001001011110100010110","0001001100010101011000","1001001100110101011000","0001001101010100011010","1001001101110100011010","0001001110010100011100","1001001110110100011100","0001001111110101110100","1001001111010100001010","0001010000110101101100","1001010000010100010010","0001010001010101100010","1001010001110101100010","0001010010010101100100","1001010010110101100100","0001010011010100100110","1001010011110100100110","0001010100010101101000","1001010100110101101000","0001010101010100101010","1001010101110100101010","0001010110010100101100","1001010110110100101100","0001010111110100101110","1001010111010101010000","0001011000110101100110","1001011000010100011000","0001011001010100110010","1001011001110100110010","0001011010010100110100","1001011010110100110100","0001011011110100110110","1001011011010101001000","0001011100010100111000","1001011100110100111000","0001011101110100111010","1001011101010101000100","0001011110110100111100","1001011110010101000010","0001011111110101101010","1001011111010100010100","0001100000111001110010","1001100000000110001100","0001100001111001011100","1001100001000110100010","0001100010111001011010","1001100010000110100100","0001100011000111000110","1001100011111001000110","0001100100111001010110","1001100100000110101000","0001100101000111001010","1001100101111001001010","0001100110000111001100","1001100110111001001100","0001100111000110001110","1001100111111001110000","0001101000111001001110","1001101000000110110000","0001101001000111010010","1001101001111001010010","0001101010000111010100","1001101010111001010100","0001101011000110010110","1001101011111000010110","0001101100000111011000","1001101100111001011000","0001101101000110011010","1001101101111000011010","0001101110000110011100","1001101110111000011100","0001101111111001110100","1001101111000110001010","0001110000111001101100","1001110000000110010010","0001110001000111100010","1001110001111001100010","0001110010000111100100","1001110010111001100100","0001110011000110100110","1001110011111000100110","0001110100000111101000","1001110100111001101000","0001110101000110101010","1001110101111000101010","0001110110000110101100","1001110110111000101100","0001110111111000101110","1001110111000111010000","0001111000111001100110","1001111000000110011000","0001111001000110110010","1001111001111000110010","0001111010000110110100","1001111010111000110100","0001111011111000110110","1001111011000111001000","0001111100000110111000","1001111100111000111000","0001111101111000111010","1001111101000111000100","0001111110111000111100","1001111110000111000010","0001111111111001101010","1001111111000110010100","0010000000001001110010","1010000000110110001100","0010000001001001011100","1010000001110110100010","0010000010001001011010","1010000010110110100100","0010000011110111000110","1010000011001001000110","0010000100001001010110","1010000100110110101000","0010000101110111001010","1010000101001001001010","0010000110110111001100","1010000110001001001100","0010000111110110001110","1010000111001001110000","0010001000001001001110","1010001000110110110000","0010001001110111010010","1010001001001001010010","0010001010110111010100","1010001010001001010100","0010001011110110010110","1010001011001000010110","0010001100110111011000","1010001100001001011000","0010001101110110011010","1010001101001000011010","0010001110110110011100","1010001110001000011100","0010001111001001110100","1010001111110110001010","0010010000001001101100","1010010000110110010010","0010010001110111100010","1010010001001001100010","0010010010110111100100","1010010010001001100100","0010010011110110100110","1010010011001000100110","0010010100110111101000","1010010100001001101000","0010010101110110101010","1010010101001000101010","0010010110110110101100","1010010110001000101100","0010010111001000101110","1010010111110111010000","0010011000001001100110","1010011000110110011000","0010011001110110110010","1010011001001000110010","0010011010110110110100","1010011010001000110100","0010011011001000110110","1010011011110111001000","0010011100110110111000","1010011100001000111000","0010011101001000111010","1010011101110111000100","0010011110001000111100","1010011110110111000010","0010011111001001101010","1010011111110110010100","0010100000101011110010","1010100000001010001100","0010100001101011011100","1010100001001010100010","0010100010101011011010","1010100010001010100100","0010100011001011000110","1010100011101011000110","0010100100101011010110","1010100100001010101000","0010100101001011001010","1010100101101011001010","0010100110001011001100","1010100110101011001100","0010100111001010001110","1010100111101011110000","0010101000101011001110","1010101000001010110000","0010101001001011010010","1010101001101011010010","0010101010001011010100","1010101010101011010100","0010101011001010010110","1010101011101010010110","0010101100001011011000","1010101100101011011000","0010101101001010011010","1010101101101010011010","0010101110001010011100","1010101110101010011100","0010101111101011110100","1010101111001010001010","0010110000101011101100","1010110000001010010010","0010110001001011100010","1010110001101011100010","0010110010001011100100","1010110010101011100100","0010110011001010100110","1010110011101010100110","0010110100001011101000","1010110100101011101000","0010110101001010101010","1010110101101010101010","0010110110001010101100","1010110110101010101100","0010110111101010101110","1010110111001011010000","0010111000101011100110","1010111000001010011000","0010111001001010110010","1010111001101010110010","0010111010001010110100","1010111010101010110100","0010111011101010110110","1010111011001011001000","0010111100001010111000","1010111100101010111000","0010111101101010111010","1010111101001011000100","0010111110101010111100","1010111110001011000010","0010111111101011101010","1010111111001010010100","0011000000101101110010","1011000000001100001100","0011000001101101011100","1011000001001100100010","0011000010101101011010","1011000010001100100100","0011000011001101000110","1011000011101101000110","0011000100101101010110","1011000100001100101000","0011000101001101001010","1011000101101101001010","0011000110001101001100","1011000110101101001100","0011000111001100001110","1011000111101101110000","0011001000101101001110","1011001000001100110000","0011001001001101010010","1011001001101101010010","0011001010001101010100","1011001010101101010100","0011001011001100010110","1011001011101100010110","0011001100001101011000","1011001100101101011000","0011001101001100011010","1011001101101100011010","0011001110001100011100","1011001110101100011100","0011001111101101110100","1011001111001100001010","0011010000101101101100","1011010000001100010010","0011010001001101100010","1011010001101101100010","0011010010001101100100","1011010010101101100100","0011010011001100100110","1011010011101100100110","0011010100001101101000","1011010100101101101000","0011010101001100101010","1011010101101100101010","0011010110001100101100","1011010110101100101100","0011010111101100101110","1011010111001101010000","0011011000101101100110","1011011000001100011000","0011011001001100110010","1011011001101100110010","0011011010001100110100","1011011010101100110100","0011011011101100110110","1011011011001101001000","0011011100001100111000","1011011100101100111000","0011011101101100111010","1011011101001101000100","0011011110101100111100","1011011110001101000010","0011011111101101101010","1011011111001100010100","0011100000010001110010","1011100000101110001100","0011100001010001011100","1011100001101110100010","0011100010010001011010","1011100010101110100100","0011100011101111000110","1011100011010001000110","0011100100010001010110","1011100100101110101000","0011100101101111001010","1011100101010001001010","0011100110101111001100","1011100110010001001100","0011100111101110001110","1011100111010001110000","0011101000010001001110","1011101000101110110000","0011101001101111010010","1011101001010001010010","0011101010101111010100","1011101010010001010100","0011101011101110010110","1011101011000010010110","0011101100101111011000","1011101100010001011000","0011101101101110011010","1011101101000010011010","0011101110101110011100","1011101110000010011100","0011101111010001110100","1011101111101110001010","0011110000010001101100","1011110000101110010010","0011110001111101100010","1011110001010001100010","0011110010111101100100","1011110010010001100100","0011110011101110100110","1011110011010000100110","0011110100111101101000","1011110100010001101000","0011110101101110101010","1011110101010000101010","0011110110101110101100","1011110110010000101100","0011110111010000101110","1011110111101111010000","0011111000010001100110","1011111000101110011000","0011111001101110110010","1011111001010000110010","0011111010101110110100","1011111010010000110100","0011111011010000110110","1011111011101111001000","0011111100101110111000","1011111100010000111000","0011111101010000111010","1011111101101111000100","0011111110010000111100","1011111110101111000010","0011111111010001101010","1011111111101110010100","0100000000000101110011","1100000000111010001101","0100000001000101011101","1100000001111010100011","0100000010000101011011","1100000010111010100101","0100000011111011000111","1100000011000101000111","0100000100000101010111","1100000100111010101001","0100000101111011001011","1100000101000101001011","0100000110111011001101","1100000110000101001101","0100000111111010001111","1100000111000101110001","0100001000000101001111","1100001000111010110001","0100001001111011010011","1100001001000101010011","0100001010111011010101","1100001010000101010101","0100001011111010010111","1100001011000100010111","0100001100111011011001","1100001100000101011001","0100001101111010011011","1100001101000100011011","0100001110111010011101","1100001110000100011101","0100001111000101110101","1100001111111010001011","0100010000000101101101","1100010000111010010011","0100010001111011100011","1100010001000101100011","0100010010111011100101","1100010010000101100101","0100010011111010100111","1100010011000100100111","0100010100111011101001","1100010100000101101001","0100010101111010101011","1100010101000100101011","0100010110111010101101","1100010110000100101101","0100010111000100101111","1100010111111011010001","0100011000000101100111","1100011000111010011001","0100011001111010110011","1100011001000100110011","0100011010111010110101","1100011010000100110101","0100011011000100110111","1100011011111011001001","0100011100000101111000","1100011100111010000110","0100011101000100111011","1100011101111011000101","0100011110000100111101","1100011110111011000011","0100011111000101101011","1100011111111010010101","0100100000110011110011","1100100000010010001101","0100100001110011011101","1100100001010010100011","0100100010110011011011","1100100010010010100101","0100100011010011000111","1100100011110011000111","0100100100110011010111","1100100100010010101001","0100100101010011001011","1100100101110011001011","0100100110010011001101","1100100110110011001101","0100100111010010001111","1100100111110011110001","0100101000110011001111","1100101000010010110001","0100101001010011010011","1100101001110011010011","0100101010010011010101","1100101010110011010101","0100101011010010010111","1100101011110010010111","0100101100010011011001","1100101100110011011001","0100101101010010011011","1100101101110010011011","0100101110010010011101","1100101110110010011101","0100101111110011110101","1100101111010010001011","0100110000110011101101","1100110000010010010011","0100110001010011100011","1100110001110011100011","0100110010010011100101","1100110010110011100101","0100110011010010100111","1100110011110010100111","0100110100010011101001","1100110100110011101001","0100110101010010101011","1100110101110010101011","0100110110010010101101","1100110110110010101101","0100110111110010101111","1100110111010011010001","0100111000110011100111","1100111000010010011001","0100111001010010110011","1100111001110010110011","0100111010010010110101","1100111010110010110101","0100111011110010110111","1100111011010011001001","0100111100110011111000","1100111100001100000110","0100111101110010111011","1100111101010011000101","0100111110110010111101","1100111110010011000011","0100111111110011101011","1100111111010010010101","0101000000110101110011","1101000000010100001101","0101000001110101011101","1101000001010100100011","0101000010110101011011","1101000010010100100101","0101000011010101000111","1101000011110101000111","0101000100110101010111","1101000100010100101001","0101000101010101001011","1101000101110101001011","0101000110010101001101","1101000110110101001101","0101000111010100001111","1101000111110101110001","0101001000110101001111","1101001000010100110001","0101001001010101010011","1101001001110101010011","0101001010010101010101","1101001010110101010101","0101001011010100010111","1101001011110100010111","0101001100010101011001","1101001100110101011001","0101001101010100011011","1101001101110100011011","0101001110010100011101","1101001110110100011101","0101001111110101110101","1101001111010100001011","0101010000110101101101","1101010000010100010011","0101010001010101100011","1101010001110101100011","0101010010010101100101","1101010010110101100101","0101010011010100100111","1101010011110100100111","0101010100010101101001","1101010100110101101001","0101010101010100101011","1101010101110100101011","0101010110010100101101","1101010110110100101101","0101010111110100101111","1101010111010101010001","0101011000110101100111","1101011000010100011001","0101011001010100110011","1101011001110100110011","0101011010010100110101","1101011010110100110101","0101011011110100110111","1101011011010101001001","0101011100110101111000","1101011100001010000110","0101011101110100111011","1101011101010101000101","0101011110110100111101","1101011110010101000011","0101011111110101101011","1101011111010100010101","0101100000111001110011","1101100000000110001101","0101100001111001011101","1101100001000110100011","0101100010111001011011","1101100010000110100101","0101100011000111000111","1101100011111001000111","0101100100111001010111","1101100100000110101001","0101100101000111001011","1101100101111001001011","0101100110000111001101","1101100110111001001101","0101100111000110001111","1101100111111001110001","0101101000111001001111","1101101000000110110001","0101101001000111010011","1101101001111001010011","0101101010000111010101","1101101010111001010101","0101101011000110010111","1101101011111000010111","0101101100000111011001","1101101100111001011001","0101101101000110011011","1101101101111000011011","0101101110000110011101","1101101110111000011101","0101101111111001110101","1101101111000110001011","0101110000111001101101","1101110000000110010011","0101110001000111100011","1101110001111001100011","0101110010000111100101","1101110010111001100101","0101110011000110100111","1101110011111000100111","0101110100000111101001","1101110100111001101001","0101110101000110101011","1101110101111000101011","0101110110000110101101","1101110110111000101101","0101110111111000101111","1101110111000111010001","0101111000111001100111","1101111000000110011001","0101111001000110110011","1101111001111000110011","0101111010000110110101","1101111010111000110101","0101111011111000110111","1101111011000111001001","0101111100111001111000","1101111100000110000110","0101111101111000111011","1101111101000111000101","0101111110111000111101","1101111110000111000011","0101111111111001101011","1101111111000110010101","0110000000001001110011","1110000000110110001101","0110000001001001011101","1110000001110110100011","0110000010001001011011","1110000010110110100101","0110000011110111000111","1110000011001001000111","0110000100001001010111","1110000100110110101001","0110000101110111001011","1110000101001001001011","0110000110110111001101","1110000110001001001101","0110000111110110001111","1110000111001001110001","0110001000001001001111","1110001000110110110001","0110001001110111010011","1110001001001001010011","0110001010110111010101","1110001010001001010101","0110001011110110010111","1110001011001000010111","0110001100110111011001","1110001100001001011001","0110001101110110011011","1110001101001000011011","0110001110110110011101","1110001110001000011101","0110001111001001110101","1110001111110110001011","0110010000001001101101","1110010000110110010011","0110010001110111100011","1110010001001001100011","0110010010110111100101","1110010010001001100101","0110010011110110100111","1110010011001000100111","0110010100110111101001","1110010100001001101001","0110010101110110101011","1110010101001000101011","0110010110110110101101","1110010110001000101101","0110010111001000101111","1110010111110111010001","0110011000001001100111","1110011000110110011001","0110011001110110110011","1110011001001000110011","0110011010110110110101","1110011010001000110101","0110011011001000110111","1110011011110111001001","0110011100001001111000","1110011100110110000110","0110011101001000111011","1110011101110111000101","0110011110001000111101","1110011110110111000011","0110011111001001101011","1110011111110110010101","0110100000101011110011","1110100000001010001101","0110100001101011011101","1110100001001010100011","0110100010101011011011","1110100010001010100101","0110100011001011000111","1110100011101011000111","0110100100101011010111","1110100100001010101001","0110100101001011001011","1110100101101011001011","0110100110001011001101","1110100110101011001101","0110100111001010001111","1110100111101011110001","0110101000101011001111","1110101000001010110001","0110101001001011010011","1110101001101011010011","0110101010001011010101","1110101010101011010101","0110101011001010010111","1110101011101010010111","0110101100001011011001","1110101100101011011001","0110101101001010011011","1110101101101010011011","0110101110001010011101","1110101110101010011101","0110101111101011110101","1110101111001010001011","0110110000101011101101","1110110000001010010011","0110110001001011100011","1110110001101011100011","0110110010001011100101","1110110010101011100101","0110110011001010100111","1110110011101010100111","0110110100001011101001","1110110100101011101001","0110110101001010101011","1110110101101010101011","0110110110001010101101","1110110110101010101101","0110110111101010101111","1110110111001011010001","0110111000101011100111","1110111000001010011001","0110111001001010110011","1110111001101010110011","0110111010001010110101","1110111010101010110101","0110111011101010110111","1110111011001011001001","0110111100101011111000","1110111100010100000110","0110111101101010111011","1110111101001011000101","0110111110101010111101","1110111110001011000011","0110111111101011101011","1110111111001010010101","0111000000101101110011","1111000000001100001101","0111000001101101011101","1111000001001100100011","0111000010101101011011","1111000010001100100101","0111000011001101000111","1111000011101101000111","0111000100101101010111","1111000100001100101001","0111000101001101001011","1111000101101101001011","0111000110001101001101","1111000110101101001101","0111000111001100001111","1111000111101101110001","0111001000101101001111","1111001000001100110001","0111001001001101010011","1111001001101101010011","0111001010001101010101","1111001010101101010101","0111001011001100010111","1111001011101100010111","0111001100001101011001","1111001100101101011001","0111001101001100011011","1111001101101100011011","0111001110001100011101","1111001110101100011101","0111001111101101110101","1111001111001100001011","0111010000101101101101","1111010000001100010011","0111010001001101100011","1111010001101101100011","0111010010001101100101","1111010010101101100101","0111010011001100100111","1111010011101100100111","0111010100001101101001","1111010100101101101001","0111010101001100101011","1111010101101100101011","0111010110001100101101","1111010110101100101101","0111010111101100101111","1111010111001101010001","0111011000101101100111","1111011000001100011001","0111011001001100110011","1111011001101100110011","0111011010001100110101","1111011010101100110101","0111011011101100110111","1111011011001101001001","0111011100101101111000","1111011100010010000110","0111011101101100111011","1111011101001101000101","0111011110101100111101","1111011110001101000011","0111011111101101101011","1111011111001100010101","0111100000010001110011","1111100000101110001101","0111100001010001011101","1111100001101110100011","0111100010010001011011","1111100010101110100101","0111100011101111000111","1111100011010001000111","0111100100010001010111","1111100100101110101001","0111100101101111001011","1111100101010001001011","0111100110101111001101","1111100110010001001101","0111100111101110001111","1111100111010001110001","0111101000010001001111","1111101000101110110001","0111101001101111010011","1111101001010001010011","0111101010101111010101","1111101010010001010101","0111101011101110010111","1111101011000010010111","0111101100101111011001","1111101100010001011001","0111101101101110011011","1111101101000010011011","0111101110101110011101","1111101110000010011101","0111101111010001110101","1111101111101110001011","0111110000010001101101","1111110000101110010011","0111110001111101100011","1111110001010001100011","0111110010111101100101","1111110010010001100101","0111110011101110100111","1111110011010000100111","0111110100111101101001","1111110100010001101001","0111110101101110101011","1111110101010000101011","0111110110101110101101","1111110110010000101101","0111110111000010101110","1111110111111101010000","0111111000010001100111","1111111000101110011001","0111111001101110110011","1111111001010000110011","0111111010101110110101","1111111010010000110101","0111111011000010110110","1111111011111101001000","0111111100000011111000","1111111100111100000110","0111111101000010111010","1111111101111101000100","0111111110000010111100","1111111110111101000010","0111111111010001101011","1111111111101110010101",
        others => (others => 'X')
    );
    type data_dec_t is array (natural range <>) of std_logic_vector(0 to 22);
    signal data_dec : data_dec_t(0 to 2047) := (
        -- dispin, d10, dispout, k, d8, err, disperr
        "0000000000000XXXXXXXX11","1000000000000XXXXXXXX11","0000000000100XXXXXXXX11","1000000000100XXXXXXXX11","0000000001000XXXXXXXX11","1000000001000XXXXXXXX11","0000000001100XXXXXXXX11","1000000001100XXXXXXXX11","0000000010000XXXXXXXX11","1000000010000XXXXXXXX11","0000000010100XXXXXXXX11","1000000010100XXXXXXXX11","0000000011000XXXXXXXX11","1000000011000XXXXXXXX11","0000000011100XXXXXXXX11","1000000011100XXXXXXXX11","0000000100000XXXXXXXX11","1000000100000XXXXXXXX11","0000000100100XXXXXXXX11","1000000100100XXXXXXXX11","0000000101000XXXXXXXX11","1000000101000XXXXXXXX11","0000000101100XXXXXXXX11","1000000101100XXXXXXXX11","0000000110000XXXXXXXX11","1000000110000XXXXXXXX11","0000000110100XXXXXXXX11","1000000110100XXXXXXXX11","0000000111000XXXXXXXX11","1000000111000XXXXXXXX11","0000000111100XXXXXXXX11","1000000111100XXXXXXXX11","0000001000000XXXXXXXX11","1000001000000XXXXXXXX11","0000001000100XXXXXXXX11","1000001000100XXXXXXXX11","0000001001000XXXXXXXX11","1000001001000XXXXXXXX11","0000001001100XXXXXXXX11","1000001001100XXXXXXXX11","0000001010000XXXXXXXX11","1000001010000XXXXXXXX11","0000001010100XXXXXXXX11","1000001010100XXXXXXXX11","0000001011000XXXXXXXX11","1000001011000XXXXXXXX11","0000001011100XXXXXXXX11","1000001011100XXXXXXXX11","0000001100000XXXXXXXX11","1000001100000XXXXXXXX11","0000001100100XXXXXXXX11","1000001100100XXXXXXXX11","0000001101000XXXXXXXX11","1000001101000XXXXXXXX11","0000001101100XXXXXXXX11","1000001101100XXXXXXXX11","0000001110000XXXXXXXX11","1000001110000XXXXXXXX11","0000001110100XXXXXXXX11","1000001110100XXXXXXXX11","0000001111000XXXXXXXX11","1000001111000XXXXXXXX11","0000001111100XXXXXXXX11","1000001111100XXXXXXXX11","0000010000000XXXXXXXX11","1000010000000XXXXXXXX11","0000010000100XXXXXXXX11","1000010000100XXXXXXXX11","0000010001000XXXXXXXX11","1000010001000XXXXXXXX11","0000010001100XXXXXXXX11","1000010001100XXXXXXXX11","0000010010000XXXXXXXX11","1000010010000XXXXXXXX11","0000010010100XXXXXXXX11","1000010010100XXXXXXXX11","0000010011000XXXXXXXX11","1000010011000XXXXXXXX11","0000010011100XXXXXXXX11","1000010011100XXXXXXXX11","0000010100000XXXXXXXX11","1000010100000XXXXXXXX11","0000010100100XXXXXXXX11","1000010100100XXXXXXXX11","0000010101000XXXXXXXX11","1000010101000XXXXXXXX11","0000010101100XXXXXXXX11","1000010101100XXXXXXXX11","0000010110000XXXXXXXX11","1000010110000XXXXXXXX11","0000010110100XXXXXXXX11","1000010110100XXXXXXXX11","0000010111000XXXXXXXX11","1000010111000XXXXXXXX11","0000010111100XXXXXXXX11","1000010111100XXXXXXXX11","0000011000000XXXXXXXX11","1000011000000XXXXXXXX11","0000011000100XXXXXXXX11","1000011000100XXXXXXXX11","0000011001000XXXXXXXX11","1000011001000XXXXXXXX11","0000011001100XXXXXXXX11","1000011001100XXXXXXXX11","0000011010000XXXXXXXX11","1000011010000XXXXXXXX11","0000011010100XXXXXXXX11","1000011010100XXXXXXXX11","0000011011000XXXXXXXX11","1000011011000XXXXXXXX11","0000011011100XXXXXXXX11","1000011011100XXXXXXXX11","0000011100000XXXXXXXX11","1000011100000XXXXXXXX11","0000011100100XXXXXXXX11","1000011100100XXXXXXXX11","0000011101000XXXXXXXX11","1000011101000XXXXXXXX11","0000011101100XXXXXXXX11","1000011101100XXXXXXXX11","0000011110000XXXXXXXX11","1000011110000XXXXXXXX11","0000011110100XXXXXXXX11","1000011110100XXXXXXXX11","0000011111000XXXXXXXX11","1000011111000XXXXXXXX11","0000011111100XXXXXXXX11","1000011111100XXXXXXXX11","0000100000000XXXXXXXX11","1000100000000XXXXXXXX11","0000100000100XXXXXXXX11","1000100000100XXXXXXXX11","0000100001000XXXXXXXX11","1000100001000XXXXXXXX11","0000100001100XXXXXXXX11","1000100001100XXXXXXXX11","0000100010000XXXXXXXX11","1000100010000XXXXXXXX11","0000100010100XXXXXXXX11","1000100010100XXXXXXXX11","0000100011000XXXXXXXX11","1000100011000XXXXXXXX11","0000100011100XXXXXXXX11","1000100011100XXXXXXXX10","0000100100000XXXXXXXX11","1000100100000XXXXXXXX11","0000100100100XXXXXXXX11","1000100100100XXXXXXXX11","0000100101000XXXXXXXX11","1000100101000XXXXXXXX11","00001001011001110101101","10001001011001110101100","0000100110000XXXXXXXX11","1000100110000XXXXXXXX11","00001001101001110110101","10001001101001110110100","00001001110001110111001","10001001110001110111000","0000100111100XXXXXXXX10","1000100111100XXXXXXXX11","0000101000000XXXXXXXX11","1000101000000XXXXXXXX11","0000101000100XXXXXXXX11","1000101000100XXXXXXXX11","0000101001000XXXXXXXX11","1000101001000XXXXXXXX11","0000101001100XXXXXXXX11","1000101001100XXXXXXXX10","0000101010000XXXXXXXX11","1000101010000XXXXXXXX11","0000101010100XXXXXXXX11","1000101010100XXXXXXXX10","0000101011000XXXXXXXX11","1000101011000XXXXXXXX10","00001010111011111011100","10001010111011111011101","0000101100000XXXXXXXX11","1000101100000XXXXXXXX11","0000101100100XXXXXXXX11","1000101100100XXXXXXXX10","0000101101000XXXXXXXX11","1000101101000XXXXXXXX10","00001011011011111101100","10001011011011111101101","0000101110000XXXXXXXX11","1000101110000XXXXXXXX10","00001011101011111110100","10001011101011111110101","00001011110011111111000","10001011110011111111001","0000101111100XXXXXXXX11","1000101111100XXXXXXXX11","0000110000000XXXXXXXX11","1000110000000XXXXXXXX11","0000110000100XXXXXXXX11","1000110000100XXXXXXXX11","0000110001000XXXXXXXX11","1000110001000XXXXXXXX11","0000110001100XXXXXXXX11","1000110001100XXXXXXXX10","0000110010000XXXXXXXX11","1000110010000XXXXXXXX11","0000110010100XXXXXXXX11","1000110010100XXXXXXXX10","0000110011000XXXXXXXX11","1000110011000XXXXXXXX10","0000110011100XXXXXXXX10","1000110011100XXXXXXXX11","0000110100000XXXXXXXX11","1000110100000XXXXXXXX11","0000110100100XXXXXXXX11","1000110100100XXXXXXXX10","0000110101000XXXXXXXX11","1000110101000XXXXXXXX10","0000110101100XXXXXXXX10","1000110101100XXXXXXXX11","0000110110000XXXXXXXX11","1000110110000XXXXXXXX10","0000110110100XXXXXXXX10","1000110110100XXXXXXXX11","0000110111000XXXXXXXX10","1000110111000XXXXXXXX11","0000110111100XXXXXXXX11","1000110111100XXXXXXXX11","0000111000000XXXXXXXX11","1000111000000XXXXXXXX11","0000111000100XXXXXXXX11","1000111000100XXXXXXXX10","0000111001000XXXXXXXX11","1000111001000XXXXXXXX10","0000111001100XXXXXXXX10","1000111001100XXXXXXXX11","0000111010000XXXXXXXX11","1000111010000XXXXXXXX10","0000111010100XXXXXXXX10","1000111010100XXXXXXXX11","0000111011000XXXXXXXX10","1000111011000XXXXXXXX11","0000111011100XXXXXXXX11","1000111011100XXXXXXXX11","0000111100000XXXXXXXX11","1000111100000XXXXXXXX10","0000111100100XXXXXXXX10","1000111100100XXXXXXXX11","0000111101000XXXXXXXX10","1000111101000XXXXXXXX11","0000111101100XXXXXXXX11","1000111101100XXXXXXXX11","00001111100011111110000","10001111100011111110001","0000111110100XXXXXXXX11","1000111110100XXXXXXXX11","0000111111000XXXXXXXX11","1000111111000XXXXXXXX11","0000111111100XXXXXXXX11","1000111111100XXXXXXXX11","0001000000000XXXXXXXX11","1001000000000XXXXXXXX11","0001000000100XXXXXXXX11","1001000000100XXXXXXXX11","0001000001000XXXXXXXX11","1001000001000XXXXXXXX11","0001000001100XXXXXXXX11","1001000001100XXXXXXXX11","0001000010000XXXXXXXX11","1001000010000XXXXXXXX11","0001000010100XXXXXXXX11","1001000010100XXXXXXXX11","0001000011000XXXXXXXX11","1001000011000XXXXXXXX11","0001000011100XXXXXXXX11","1001000011100XXXXXXXX10","0001000100000XXXXXXXX11","1001000100000XXXXXXXX11","0001000100100XXXXXXXX11","1001000100100XXXXXXXX11","0001000101000XXXXXXXX11","1001000101000XXXXXXXX11","00010001011000000101101","10010001011000000101100","0001000110000XXXXXXXX11","1001000110000XXXXXXXX11","00010001101000000110101","10010001101000000110100","00010001110000000111001","10010001110000000111000","0001000111100XXXXXXXX10","1001000111100XXXXXXXX11","0001001000000XXXXXXXX11","1001001000000XXXXXXXX11","0001001000100XXXXXXXX11","1001001000100XXXXXXXX11","0001001001000XXXXXXXX11","1001001001000XXXXXXXX11","00010010011000001001101","10010010011000001001100","0001001010000XXXXXXXX11","1001001010000XXXXXXXX11","00010010101000001010101","10010010101000001010100","00010010110000001011001","10010010110000001011000","00010010111000001011100","10010010111000001011101","0001001100000XXXXXXXX11","1001001100000XXXXXXXX11","00010011001000001100101","10010011001000001100100","00010011010000001101001","10010011010000001101000","00010011011000001101100","10010011011000001101101","00010011100000001110001","10010011100000001110000","00010011101000001110100","10010011101000001110101","00010011110000001111000","10010011110000001111001","0001001111100XXXXXXXX11","1001001111100XXXXXXXX11","0001010000000XXXXXXXX11","1001010000000XXXXXXXX11","0001010000100XXXXXXXX11","1001010000100XXXXXXXX11","0001010001000XXXXXXXX11","1001010001000XXXXXXXX11","00010100011000000001101","10010100011000000001100","0001010010000XXXXXXXX11","1001010010000XXXXXXXX11","00010100101000000010101","10010100101000000010100","00010100110000000011001","10010100110000000011000","00010100111000000100000","10010100111000000100001","0001010100000XXXXXXXX11","1001010100000XXXXXXXX11","00010101001000000100101","10010101001000000100100","00010101010000000101001","10010101010000000101000","00010101011000000010000","10010101011000000010001","00010101100000000110001","10010101100000000110000","00010101101000000001000","10010101101000000001001","00010101110000000000100","10010101110000000000101","0001010111100XXXXXXXX11","1001010111100XXXXXXXX11","0001011000000XXXXXXXX11","1001011000000XXXXXXXX11","00010110001000001000101","10010110001000001000100","00010110010000001001001","10010110010000001001000","00010110011000001100000","10010110011000001100001","00010110100000001010001","10010110100000001010000","00010110101000001111100","10010110101000001111101","00010110110000001000000","10010110110000001000001","0001011011100XXXXXXXX11","1001011011100XXXXXXXX11","00010111000000000011101","10010111000000000011100","00010111001000000000000","10010111001000000000001","00010111010000000111100","10010111010000000111101","0001011101100XXXXXXXX11","1001011101100XXXXXXXX11","00010111100010001110000","10010111100010001110001","0001011110100XXXXXXXX11","1001011110100XXXXXXXX11","0001011111000XXXXXXXX11","1001011111000XXXXXXXX11","0001011111100XXXXXXXX11","1001011111100XXXXXXXX11","0001100000000XXXXXXXX11","1001100000000XXXXXXXX11","0001100000100XXXXXXXX11","1001100000100XXXXXXXX11","0001100001000XXXXXXXX11","1001100001000XXXXXXXX11","00011000011010111110001","10011000011010111110000","0001100010000XXXXXXXX11","1001100010000XXXXXXXX11","00011000101000110111101","10011000101000110111100","00011000110000110000001","10011000110000110000000","00011000111000110011100","10011000111100110011101","0001100100000XXXXXXXX11","1001100100000XXXXXXXX11","00011001001000111000001","10011001001000111000000","00011001010000111111101","10011001010000111111100","00011001011000110101100","10011001011100110101101","00011001100000111100001","10011001100000111100000","00011001101000110110100","10011001101100110110101","00011001110000110111000","10011001110100110111001","0001100111110XXXXXXXX10","1001100111110XXXXXXXX11","0001101000000XXXXXXXX11","1001101000000XXXXXXXX11","00011010001000110000101","10011010001000110000100","00011010010000110001001","10011010010000110001000","00011010011000111001100","10011010011100111001101","00011010100000110010001","10011010100000110010000","00011010101000111010100","10011010101100111010101","00011010110000111011000","10011010110100111011001","0001101011110XXXXXXXX10","1001101011110XXXXXXXX11","00011011000000110100001","10011011000000110100000","00011011001000111100100","10011011001100111100101","00011011010000111101000","10011011010100111101001","0001101101110XXXXXXXX10","1001101101110XXXXXXXX11","00011011100000111110000","10011011100100111110001","0001101110110XXXXXXXX10","1001101110110XXXXXXXX11","0001101111010XXXXXXXX10","1001101111010XXXXXXXX11","0001101111110XXXXXXXX11","1001101111110XXXXXXXX11","0001110000000XXXXXXXX11","1001110000000XXXXXXXX11","00011100001000111111001","10011100001000111111000","00011100010000111110101","10011100010000111110100","00011100011000110001100","10011100011100110001101","00011100100000111101101","10011100100000111101100","00011100101000110010100","10011100101100110010101","00011100110000110011000","10011100110100110011001","0001110011110XXXXXXXX10","1001110011110XXXXXXXX11","00011101000000111011101","10011101000000111011100","00011101001000110100100","10011101001100110100101","00011101010000110101000","10011101010100110101001","0001110101110XXXXXXXX10","1001110101110XXXXXXXX11","00011101100000110110000","10011101100100110110001","0001110110110XXXXXXXX10","1001110110110XXXXXXXX11","0001110111010XXXXXXXX10","1001110111010XXXXXXXX11","0001110111110XXXXXXXX11","1001110111110XXXXXXXX11","0001111000000XXXXXXXX11","1001111000000XXXXXXXX10","00011110001000111000100","10011110001100111000101","00011110010000111001000","10011110010100111001001","0001111001110XXXXXXXX10","1001111001110XXXXXXXX11","00011110100000111010000","10011110100100111010001","0001111010110XXXXXXXX10","1001111010110XXXXXXXX11","0001111011010XXXXXXXX10","1001111011010XXXXXXXX11","0001111011110XXXXXXXX11","1001111011110XXXXXXXX11","0001111100000XXXXXXXX10","1001111100010XXXXXXXX10","0001111100110XXXXXXXX10","1001111100110XXXXXXXX11","0001111101010XXXXXXXX10","1001111101010XXXXXXXX11","0001111101110XXXXXXXX11","1001111101110XXXXXXXX11","0001111110010XXXXXXXX10","1001111110010XXXXXXXX11","0001111110110XXXXXXXX11","1001111110110XXXXXXXX11","0001111111010XXXXXXXX11","1001111111010XXXXXXXX11","0001111111110XXXXXXXX11","1001111111110XXXXXXXX11","0010000000000XXXXXXXX11","1010000000000XXXXXXXX11","0010000000100XXXXXXXX11","1010000000100XXXXXXXX11","0010000001000XXXXXXXX11","1010000001000XXXXXXXX11","0010000001100XXXXXXXX11","1010000001100XXXXXXXX11","0010000010000XXXXXXXX11","1010000010000XXXXXXXX11","0010000010100XXXXXXXX11","1010000010100XXXXXXXX11","0010000011000XXXXXXXX11","1010000011000XXXXXXXX11","0010000011100XXXXXXXX11","1010000011100XXXXXXXX10","0010000100000XXXXXXXX11","1010000100000XXXXXXXX11","0010000100100XXXXXXXX11","1010000100100XXXXXXXX11","0010000101000XXXXXXXX11","1010000101000XXXXXXXX11","00100001011001000101101","10100001011001000101100","0010000110000XXXXXXXX11","1010000110000XXXXXXXX11","00100001101001000110101","10100001101001000110100","00100001110001000111001","10100001110001000111000","0010000111100XXXXXXXX10","1010000111100XXXXXXXX11","0010001000000XXXXXXXX11","1010001000000XXXXXXXX11","0010001000100XXXXXXXX11","1010001000100XXXXXXXX11","0010001001000XXXXXXXX11","1010001001000XXXXXXXX11","00100010011001001001101","10100010011001001001100","0010001010000XXXXXXXX11","1010001010000XXXXXXXX11","00100010101001001010101","10100010101001001010100","00100010110001001011001","10100010110001001011000","00100010111001001011100","10100010111001001011101","0010001100000XXXXXXXX11","1010001100000XXXXXXXX11","00100011001001001100101","10100011001001001100100","00100011010001001101001","10100011010001001101000","00100011011001001101100","10100011011001001101101","00100011100001001110001","10100011100001001110000","00100011101001001110100","10100011101001001110101","00100011110001001111000","10100011110001001111001","0010001111100XXXXXXXX11","1010001111100XXXXXXXX11","0010010000000XXXXXXXX11","1010010000000XXXXXXXX11","0010010000100XXXXXXXX11","1010010000100XXXXXXXX11","0010010001000XXXXXXXX11","1010010001000XXXXXXXX11","00100100011001000001101","10100100011001000001100","0010010010000XXXXXXXX11","1010010010000XXXXXXXX11","00100100101001000010101","10100100101001000010100","00100100110001000011001","10100100110001000011000","00100100111001000100000","10100100111001000100001","0010010100000XXXXXXXX11","1010010100000XXXXXXXX11","00100101001001000100101","10100101001001000100100","00100101010001000101001","10100101010001000101000","00100101011001000010000","10100101011001000010001","00100101100001000110001","10100101100001000110000","00100101101001000001000","10100101101001000001001","00100101110001000000100","10100101110001000000101","0010010111100XXXXXXXX11","1010010111100XXXXXXXX11","0010011000000XXXXXXXX11","1010011000000XXXXXXXX11","00100110001001001000101","10100110001001001000100","00100110010001001001001","10100110010001001001000","00100110011001001100000","10100110011001001100001","00100110100001001010001","10100110100001001010000","00100110101001001111100","10100110101001001111101","00100110110001001000000","10100110110001001000001","0010011011100XXXXXXXX11","1010011011100XXXXXXXX11","00100111000001000011101","10100111000001000011100","00100111001001000000000","10100111001001000000001","00100111010001000111100","10100111010001000111101","0010011101100XXXXXXXX11","1010011101100XXXXXXXX11","00100111100011001110000","10100111100011001110001","0010011110100XXXXXXXX11","1010011110100XXXXXXXX11","0010011111000XXXXXXXX11","1010011111000XXXXXXXX11","0010011111100XXXXXXXX11","1010011111100XXXXXXXX11","0010100000000XXXXXXXX11","1010100000000XXXXXXXX11","0010100000100XXXXXXXX11","1010100000100XXXXXXXX11","0010100001000XXXXXXXX11","1010100001000XXXXXXXX11","00101000011010101110001","10101000011010101110000","0010100010000XXXXXXXX11","1010100010000XXXXXXXX11","00101000101001010111101","10101000101001010111100","00101000110001010000001","10101000110001010000000","00101000111001010011100","10101000111101010011101","0010100100000XXXXXXXX11","1010100100000XXXXXXXX11","00101001001001011000001","10101001001001011000000","00101001010001011111101","10101001010001011111100","00101001011001010101100","10101001011101010101100","00101001100001011100001","10101001100001011100000","00101001101001010110100","10101001101101010110100","00101001110001010111000","10101001110101010111000","0010100111110XXXXXXXX10","1010100111110XXXXXXXX11","0010101000000XXXXXXXX11","1010101000000XXXXXXXX11","00101010001001010000101","10101010001001010000100","00101010010001010001001","10101010010001010001000","00101010011001011001100","10101010011101011001100","00101010100001010010001","10101010100001010010000","00101010101001011010100","10101010101101011010100","00101010110001011011000","10101010110101011011000","00101010111101011011100","10101010111101011011101","00101011000001010100001","10101011000001010100000","00101011001001011100100","10101011001101011100100","00101011010001011101000","10101011010101011101000","00101011011101011101100","10101011011101011101101","00101011100001011110000","10101011100101011110000","00101011101101011110100","10101011101101011110101","00101011110101011111000","10101011110101011111001","0010101111110XXXXXXXX11","1010101111110XXXXXXXX11","0010110000000XXXXXXXX11","1010110000000XXXXXXXX11","00101100001001011111001","10101100001001011111000","00101100010001011110101","10101100010001011110100","00101100011001010001100","10101100011101010001100","00101100100001011101101","10101100100001011101100","00101100101001010010100","10101100101101010010100","00101100110001010011000","10101100110101010011000","00101100111101010100000","10101100111101010100001","00101101000001011011101","10101101000001011011100","00101101001001010100100","10101101001101010100100","00101101010001010101000","10101101010101010101000","00101101011101010010000","10101101011101010010001","00101101100001010110000","10101101100101010110000","00101101101101010001000","10101101101101010001001","00101101110101010000100","10101101110101010000101","0010110111110XXXXXXXX11","1010110111110XXXXXXXX11","0010111000000XXXXXXXX11","1010111000000XXXXXXXX10","00101110001001011000100","10101110001101011000100","00101110010001011001000","10101110010101011001000","00101110011101011100000","10101110011101011100001","00101110100001011010000","10101110100101011010000","00101110101101011111100","10101110101101011111101","00101110110101011000000","10101110110101011000001","0010111011110XXXXXXXX11","1010111011110XXXXXXXX11","00101111000001010011101","10101111000101010011100","00101111001101010000000","10101111001101010000001","00101111010101010111100","10101111010101010111101","0010111101110XXXXXXXX11","1010111101110XXXXXXXX11","00101111100111011110000","10101111100111011110001","0010111110110XXXXXXXX11","1010111110110XXXXXXXX11","0010111111010XXXXXXXX11","1010111111010XXXXXXXX11","0010111111110XXXXXXXX11","1010111111110XXXXXXXX11","0011000000000XXXXXXXX11","1011000000000XXXXXXXX11","0011000000100XXXXXXXX11","1011000000100XXXXXXXX11","0011000001000XXXXXXXX11","1011000001000XXXXXXXX11","00110000011010011110001","10110000011010011110000","0011000010000XXXXXXXX11","1011000010000XXXXXXXX11","00110000101001100111101","10110000101001100111100","00110000110001100000001","10110000110001100000000","00110000111001100011100","10110000111101100011101","0011000100000XXXXXXXX11","1011000100000XXXXXXXX11","00110001001001101000001","10110001001001101000000","00110001010001101111101","10110001010001101111100","00110001011001100101100","10110001011101100101100","00110001100001101100001","10110001100001101100000","00110001101001100110100","10110001101101100110100","00110001110001100111000","10110001110101100111000","0011000111110XXXXXXXX10","1011000111110XXXXXXXX11","0011001000000XXXXXXXX11","1011001000000XXXXXXXX11","00110010001001100000101","10110010001001100000100","00110010010001100001001","10110010010001100001000","00110010011001101001100","10110010011101101001100","00110010100001100010001","10110010100001100010000","00110010101001101010100","10110010101101101010100","00110010110001101011000","10110010110101101011000","00110010111101101011100","10110010111101101011101","00110011000001100100001","10110011000001100100000","00110011001001101100100","10110011001101101100100","00110011010001101101000","10110011010101101101000","00110011011101101101100","10110011011101101101101","00110011100001101110000","10110011100101101110000","00110011101101101110100","10110011101101101110101","00110011110101101111000","10110011110101101111001","0011001111110XXXXXXXX11","1011001111110XXXXXXXX11","0011010000000XXXXXXXX11","1011010000000XXXXXXXX11","00110100001001101111001","10110100001001101111000","00110100010001101110101","10110100010001101110100","00110100011001100001100","10110100011101100001100","00110100100001101101101","10110100100001101101100","00110100101001100010100","10110100101101100010100","00110100110001100011000","10110100110101100011000","00110100111101100100000","10110100111101100100001","00110101000001101011101","10110101000001101011100","00110101001001100100100","10110101001101100100100","00110101010001100101000","10110101010101100101000","00110101011101100010000","10110101011101100010001","00110101100001100110000","10110101100101100110000","00110101101101100001000","10110101101101100001001","00110101110101100000100","10110101110101100000101","0011010111110XXXXXXXX11","1011010111110XXXXXXXX11","0011011000000XXXXXXXX11","1011011000000XXXXXXXX10","00110110001001101000100","10110110001101101000100","00110110010001101001000","10110110010101101001000","00110110011101101100000","10110110011101101100001","00110110100001101010000","10110110100101101010000","00110110101101101111100","10110110101101101111101","00110110110101101000000","10110110110101101000001","0011011011110XXXXXXXX11","1011011011110XXXXXXXX11","00110111000001100011101","10110111000101100011100","00110111001101100000000","10110111001101100000001","00110111010101100111100","10110111010101100111101","0011011101110XXXXXXXX11","1011011101110XXXXXXXX11","00110111100111101110000","10110111100111101110001","0011011110110XXXXXXXX11","1011011110110XXXXXXXX11","0011011111010XXXXXXXX11","1011011111010XXXXXXXX11","0011011111110XXXXXXXX11","1011011111110XXXXXXXX11","0011100000010XXXXXXXX11","1011100000010XXXXXXXX11","0011100000110XXXXXXXX11","1011100000110XXXXXXXX11","0011100001010XXXXXXXX11","1011100001010XXXXXXXX11","0011100001110XXXXXXXX11","1011100001110XXXXXXXX10","0011100010010XXXXXXXX11","1011100010010XXXXXXXX11","00111000101101110111101","10111000101101110111100","00111000110101110000001","10111000110101110000000","00111000111101110011100","10111000111101110011101","0011100100010XXXXXXXX11","1011100100010XXXXXXXX11","00111001001101111000001","10111001001101111000000","00111001010101111111101","10111001010101111111100","00111001011101110101100","10111001011101110101101","00111001100101111100001","10111001100101111100000","00111001101101110110100","10111001101101110110101","00111001110101110111000","10111001110101110111001","0011100111110XXXXXXXX11","1011100111110XXXXXXXX11","0011101000010XXXXXXXX11","1011101000010XXXXXXXX11","00111010001101110000101","10111010001101110000100","00111010010101110001001","10111010010101110001000","00111010011101111001100","10111010011101111001101","00111010100101110010001","10111010100101110010000","00111010101101111010100","10111010101101111010101","00111010110101111011000","10111010110101111011001","0011101011110XXXXXXXX11","1011101011110XXXXXXXX11","00111011000101110100001","10111011000101110100000","00111011001101111100100","10111011001101111100101","00111011010101111101000","10111011010101111101001","0011101101110XXXXXXXX11","1011101101110XXXXXXXX11","00111011100101111110000","10111011100101111110001","0011101110110XXXXXXXX11","1011101110110XXXXXXXX11","0011101111010XXXXXXXX11","1011101111010XXXXXXXX11","0011101111110XXXXXXXX11","1011101111110XXXXXXXX11","0011110000010XXXXXXXX11","1011110000010XXXXXXXX11","00111100001101111111001","10111100001101111111000","00111100010101111110101","10111100010101111110100","00111100011101110001100","10111100011101110001101","00111100100101111101101","10111100100101111101100","00111100101101110010100","10111100101101110010101","00111100110101110011000","10111100110101110011001","0011110011110XXXXXXXX11","1011110011110XXXXXXXX11","00111101000101111011101","10111101000101111011100","00111101001101110100100","10111101001101110100101","00111101010101110101000","10111101010101110101001","0011110101110XXXXXXXX11","1011110101110XXXXXXXX11","00111101100101110110000","10111101100101110110001","0011110110110XXXXXXXX11","1011110110110XXXXXXXX11","0011110111010XXXXXXXX11","1011110111010XXXXXXXX11","0011110111110XXXXXXXX11","1011110111110XXXXXXXX11","0011111000010XXXXXXXX11","1011111000010XXXXXXXX10","0011111000110XXXXXXXX10","1011111000110XXXXXXXX11","0011111001010XXXXXXXX10","1011111001010XXXXXXXX11","0011111001110XXXXXXXX11","1011111001110XXXXXXXX11","0011111010010XXXXXXXX10","1011111010010XXXXXXXX11","0011111010110XXXXXXXX11","1011111010110XXXXXXXX11","0011111011010XXXXXXXX11","1011111011010XXXXXXXX11","0011111011110XXXXXXXX11","1011111011110XXXXXXXX11","0011111100010XXXXXXXX10","1011111100010XXXXXXXX11","0011111100110XXXXXXXX11","1011111100110XXXXXXXX11","0011111101010XXXXXXXX11","1011111101010XXXXXXXX11","0011111101110XXXXXXXX11","1011111101110XXXXXXXX11","0011111110010XXXXXXXX11","1011111110010XXXXXXXX11","0011111110110XXXXXXXX11","1011111110110XXXXXXXX11","0011111111010XXXXXXXX11","1011111111010XXXXXXXX11","0011111111110XXXXXXXX11","1011111111110XXXXXXXX11","0100000000000XXXXXXXX11","1100000000000XXXXXXXX11","0100000000100XXXXXXXX11","1100000000100XXXXXXXX11","0100000001000XXXXXXXX11","1100000001000XXXXXXXX11","0100000001100XXXXXXXX11","1100000001100XXXXXXXX11","0100000010000XXXXXXXX11","1100000010000XXXXXXXX11","0100000010100XXXXXXXX11","1100000010100XXXXXXXX11","0100000011000XXXXXXXX11","1100000011000XXXXXXXX11","0100000011100XXXXXXXX11","1100000011100XXXXXXXX10","0100000100000XXXXXXXX11","1100000100000XXXXXXXX11","0100000100100XXXXXXXX11","1100000100100XXXXXXXX11","0100000101000XXXXXXXX11","1100000101000XXXXXXXX11","0100000101100XXXXXXXX11","1100000101100XXXXXXXX10","0100000110000XXXXXXXX11","1100000110000XXXXXXXX11","0100000110100XXXXXXXX11","1100000110100XXXXXXXX10","0100000111000XXXXXXXX11","1100000111000XXXXXXXX10","0100000111100XXXXXXXX10","1100000111100XXXXXXXX11","0100001000000XXXXXXXX11","1100001000000XXXXXXXX11","0100001000100XXXXXXXX11","1100001000100XXXXXXXX11","0100001001000XXXXXXXX11","1100001001000XXXXXXXX11","01000010011001111001101","11000010011001111001100","0100001010000XXXXXXXX11","1100001010000XXXXXXXX11","01000010101001111010101","11000010101001111010100","01000010110001111011001","11000010110001111011000","01000010111001111011100","11000010111001111011101","0100001100000XXXXXXXX11","1100001100000XXXXXXXX11","01000011001001111100101","11000011001001111100100","01000011010001111101001","11000011010001111101000","01000011011001111101100","11000011011001111101101","01000011100001111110001","11000011100001111110000","01000011101001111110100","11000011101001111110101","01000011110001111111000","11000011110001111111001","0100001111100XXXXXXXX11","1100001111100XXXXXXXX11","0100010000000XXXXXXXX11","1100010000000XXXXXXXX11","0100010000100XXXXXXXX11","1100010000100XXXXXXXX11","0100010001000XXXXXXXX11","1100010001000XXXXXXXX11","01000100011001110001101","11000100011001110001100","0100010010000XXXXXXXX11","1100010010000XXXXXXXX11","01000100101001110010101","11000100101001110010100","01000100110001110011001","11000100110001110011000","01000100111001110100000","11000100111001110100001","0100010100000XXXXXXXX11","1100010100000XXXXXXXX11","01000101001001110100101","11000101001001110100100","01000101010001110101001","11000101010001110101000","01000101011001110010000","11000101011001110010001","01000101100001110110001","11000101100001110110000","01000101101001110001000","11000101101001110001001","01000101110001110000100","11000101110001110000101","0100010111100XXXXXXXX11","1100010111100XXXXXXXX11","0100011000000XXXXXXXX11","1100011000000XXXXXXXX11","01000110001001111000101","11000110001001111000100","01000110010001111001001","11000110010001111001000","01000110011001111100000","11000110011001111100001","01000110100001111010001","11000110100001111010000","01000110101001111111100","11000110101001111111101","01000110110001111000000","11000110110001111000001","0100011011100XXXXXXXX11","1100011011100XXXXXXXX11","01000111000001110011101","11000111000001110011100","01000111001001110000000","11000111001001110000001","01000111010001110111100","11000111010001110111101","0100011101100XXXXXXXX11","1100011101100XXXXXXXX11","0100011110000XXXXXXXX10","1100011110000XXXXXXXX11","0100011110100XXXXXXXX11","1100011110100XXXXXXXX11","0100011111000XXXXXXXX11","1100011111000XXXXXXXX11","0100011111100XXXXXXXX11","1100011111100XXXXXXXX11","0100100000000XXXXXXXX11","1100100000000XXXXXXXX11","0100100000100XXXXXXXX11","1100100000100XXXXXXXX11","0100100001000XXXXXXXX11","1100100001000XXXXXXXX11","01001000011011101110001","11001000011011101110000","0100100010000XXXXXXXX11","1100100010000XXXXXXXX11","01001000101000010111101","11001000101000010111100","01001000110000010000001","11001000110000010000000","01001000111000010011100","11001000111100010011101","0100100100000XXXXXXXX11","1100100100000XXXXXXXX11","01001001001000011000001","11001001001000011000000","01001001010000011111101","11001001010000011111100","01001001011000010101100","11001001011100010101100","01001001100000011100001","11001001100000011100000","01001001101000010110100","11001001101100010110100","01001001110000010111000","11001001110100010111000","0100100111110XXXXXXXX10","1100100111110XXXXXXXX11","0100101000000XXXXXXXX11","1100101000000XXXXXXXX11","01001010001000010000101","11001010001000010000100","01001010010000010001001","11001010010000010001000","01001010011000011001100","11001010011100011001100","01001010100000010010001","11001010100000010010000","01001010101000011010100","11001010101100011010100","01001010110000011011000","11001010110100011011000","01001010111100011011100","11001010111100011011101","01001011000000010100001","11001011000000010100000","01001011001000011100100","11001011001100011100100","01001011010000011101000","11001011010100011101000","01001011011100011101100","11001011011100011101101","01001011100000011110000","11001011100100011110000","01001011101100011110100","11001011101100011110101","01001011110100011111000","11001011110100011111001","0100101111110XXXXXXXX11","1100101111110XXXXXXXX11","0100110000000XXXXXXXX11","1100110000000XXXXXXXX11","01001100001000011111001","11001100001000011111000","01001100010000011110101","11001100010000011110100","01001100011000010001100","11001100011100010001100","01001100100000011101101","11001100100000011101100","01001100101000010010100","11001100101100010010100","01001100110000010011000","11001100110100010011000","01001100111100010100000","11001100111100010100001","01001101000000011011101","11001101000000011011100","01001101001000010100100","11001101001100010100100","01001101010000010101000","11001101010100010101000","01001101011100010010000","11001101011100010010001","01001101100000010110000","11001101100100010110000","01001101101100010001000","11001101101100010001001","01001101110100010000100","11001101110100010000101","0100110111110XXXXXXXX11","1100110111110XXXXXXXX11","0100111000000XXXXXXXX11","1100111000000XXXXXXXX10","01001110001000011000100","11001110001100011000100","01001110010000011001000","11001110010100011001000","01001110011100011100000","11001110011100011100001","01001110100000011010000","11001110100100011010000","01001110101100011111100","11001110101100011111101","01001110110100011000000","11001110110100011000001","0100111011110XXXXXXXX11","1100111011110XXXXXXXX11","01001111000000010011101","11001111000100010011100","01001111001100010000000","11001111001100010000001","01001111010100010111100","11001111010100010111101","0100111101110XXXXXXXX11","1100111101110XXXXXXXX11","01001111100110011110000","11001111100110011110001","0100111110110XXXXXXXX11","1100111110110XXXXXXXX11","0100111111010XXXXXXXX11","1100111111010XXXXXXXX11","0100111111110XXXXXXXX11","1100111111110XXXXXXXX11","0101000000000XXXXXXXX11","1101000000000XXXXXXXX11","0101000000100XXXXXXXX11","1101000000100XXXXXXXX11","0101000001000XXXXXXXX11","1101000001000XXXXXXXX11","01010000011011011110001","11010000011011011110000","0101000010000XXXXXXXX11","1101000010000XXXXXXXX11","01010000101000100111101","11010000101000100111100","01010000110000100000001","11010000110000100000000","01010000111000100011100","11010000111100100011101","0101000100000XXXXXXXX11","1101000100000XXXXXXXX11","01010001001000101000001","11010001001000101000000","01010001010000101111101","11010001010000101111100","01010001011000100101100","11010001011100100101100","01010001100000101100001","11010001100000101100000","01010001101000100110100","11010001101100100110100","01010001110000100111000","11010001110100100111000","0101000111110XXXXXXXX10","1101000111110XXXXXXXX11","0101001000000XXXXXXXX11","1101001000000XXXXXXXX11","01010010001000100000101","11010010001000100000100","01010010010000100001001","11010010010000100001000","01010010011000101001100","11010010011100101001100","01010010100000100010001","11010010100000100010000","01010010101000101010100","11010010101100101010100","01010010110000101011000","11010010110100101011000","01010010111100101011100","11010010111100101011101","01010011000000100100001","11010011000000100100000","01010011001000101100100","11010011001100101100100","01010011010000101101000","11010011010100101101000","01010011011100101101100","11010011011100101101101","01010011100000101110000","11010011100100101110000","01010011101100101110100","11010011101100101110101","01010011110100101111000","11010011110100101111001","0101001111110XXXXXXXX11","1101001111110XXXXXXXX11","0101010000000XXXXXXXX11","1101010000000XXXXXXXX11","01010100001000101111001","11010100001000101111000","01010100010000101110101","11010100010000101110100","01010100011000100001100","11010100011100100001100","01010100100000101101101","11010100100000101101100","01010100101000100010100","11010100101100100010100","01010100110000100011000","11010100110100100011000","01010100111100100100000","11010100111100100100001","01010101000000101011101","11010101000000101011100","01010101001000100100100","11010101001100100100100","01010101010000100101000","11010101010100100101000","01010101011100100010000","11010101011100100010001","01010101100000100110000","11010101100100100110000","01010101101100100001000","11010101101100100001001","01010101110100100000100","11010101110100100000101","0101010111110XXXXXXXX11","1101010111110XXXXXXXX11","0101011000000XXXXXXXX11","1101011000000XXXXXXXX10","01010110001000101000100","11010110001100101000100","01010110010000101001000","11010110010100101001000","01010110011100101100000","11010110011100101100001","01010110100000101010000","11010110100100101010000","01010110101100101111100","11010110101100101111101","01010110110100101000000","11010110110100101000001","0101011011110XXXXXXXX11","1101011011110XXXXXXXX11","01010111000000100011101","11010111000100100011100","01010111001100100000000","11010111001100100000001","01010111010100100111100","11010111010100100111101","0101011101110XXXXXXXX11","1101011101110XXXXXXXX11","01010111100110101110000","11010111100110101110001","0101011110110XXXXXXXX11","1101011110110XXXXXXXX11","0101011111010XXXXXXXX11","1101011111010XXXXXXXX11","0101011111110XXXXXXXX11","1101011111110XXXXXXXX11","0101100000010XXXXXXXX11","1101100000010XXXXXXXX11","0101100000110XXXXXXXX11","1101100000110XXXXXXXX11","0101100001010XXXXXXXX11","1101100001010XXXXXXXX11","01011000011111001110001","11011000011111001110000","0101100010010XXXXXXXX11","1101100010010XXXXXXXX11","01011000101101000111101","11011000101101000111100","01011000110101000000001","11011000110101000000000","01011000111101000011100","11011000111101000011101","0101100100010XXXXXXXX11","1101100100010XXXXXXXX11","01011001001101001000001","11011001001101001000000","01011001010101001111101","11011001010101001111100","01011001011101000101100","11011001011101000101101","01011001100101001100001","11011001100101001100000","01011001101101000110100","11011001101101000110101","01011001110101000111000","11011001110101000111001","0101100111110XXXXXXXX11","1101100111110XXXXXXXX11","0101101000010XXXXXXXX11","1101101000010XXXXXXXX11","01011010001101000000101","11011010001101000000100","01011010010101000001001","11011010010101000001000","01011010011101001001100","11011010011101001001101","01011010100101000010001","11011010100101000010000","01011010101101001010100","11011010101101001010101","01011010110101001011000","11011010110101001011001","0101101011110XXXXXXXX11","1101101011110XXXXXXXX11","01011011000101000100001","11011011000101000100000","01011011001101001100100","11011011001101001100101","01011011010101001101000","11011011010101001101001","0101101101110XXXXXXXX11","1101101101110XXXXXXXX11","01011011100101001110000","11011011100101001110001","0101101110110XXXXXXXX11","1101101110110XXXXXXXX11","0101101111010XXXXXXXX11","1101101111010XXXXXXXX11","0101101111110XXXXXXXX11","1101101111110XXXXXXXX11","0101110000010XXXXXXXX11","1101110000010XXXXXXXX11","01011100001101001111001","11011100001101001111000","01011100010101001110101","11011100010101001110100","01011100011101000001100","11011100011101000001101","01011100100101001101101","11011100100101001101100","01011100101101000010100","11011100101101000010101","01011100110101000011000","11011100110101000011001","0101110011110XXXXXXXX11","1101110011110XXXXXXXX11","01011101000101001011101","11011101000101001011100","01011101001101000100100","11011101001101000100101","01011101010101000101000","11011101010101000101001","0101110101110XXXXXXXX11","1101110101110XXXXXXXX11","01011101100101000110000","11011101100101000110001","0101110110110XXXXXXXX11","1101110110110XXXXXXXX11","0101110111010XXXXXXXX11","1101110111010XXXXXXXX11","0101110111110XXXXXXXX11","1101110111110XXXXXXXX11","0101111000010XXXXXXXX11","1101111000010XXXXXXXX10","01011110001101001000100","11011110001101001000101","01011110010101001001000","11011110010101001001001","0101111001110XXXXXXXX11","1101111001110XXXXXXXX11","01011110100101001010000","11011110100101001010001","0101111010110XXXXXXXX11","1101111010110XXXXXXXX11","0101111011010XXXXXXXX11","1101111011010XXXXXXXX11","0101111011110XXXXXXXX11","1101111011110XXXXXXXX11","0101111100010XXXXXXXX10","1101111100010XXXXXXXX11","0101111100110XXXXXXXX11","1101111100110XXXXXXXX11","0101111101010XXXXXXXX11","1101111101010XXXXXXXX11","0101111101110XXXXXXXX11","1101111101110XXXXXXXX11","0101111110010XXXXXXXX11","1101111110010XXXXXXXX11","0101111110110XXXXXXXX11","1101111110110XXXXXXXX11","0101111111010XXXXXXXX11","1101111111010XXXXXXXX11","0101111111110XXXXXXXX11","1101111111110XXXXXXXX11","0110000000000XXXXXXXX11","1110000000000XXXXXXXX11","0110000000100XXXXXXXX11","1110000000100XXXXXXXX11","0110000001000XXXXXXXX11","1110000001000XXXXXXXX11","0110000001100XXXXXXXX11","1110000001100XXXXXXXX10","0110000010000XXXXXXXX11","1110000010000XXXXXXXX11","0110000010100XXXXXXXX11","1110000010100XXXXXXXX10","0110000011000XXXXXXXX11","1110000011000XXXXXXXX10","0110000011100XXXXXXXX10","1110000011110XXXXXXXX10","0110000100000XXXXXXXX11","1110000100000XXXXXXXX11","0110000100100XXXXXXXX11","1110000100100XXXXXXXX10","0110000101000XXXXXXXX11","1110000101000XXXXXXXX10","01100001011000110101101","11100001011100110101100","0110000110000XXXXXXXX11","1110000110000XXXXXXXX10","01100001101000110110101","11100001101100110110100","01100001110000110111001","11100001110100110111000","0110000111110XXXXXXXX10","1110000111110XXXXXXXX11","0110001000000XXXXXXXX11","1110001000000XXXXXXXX11","0110001000100XXXXXXXX11","1110001000100XXXXXXXX10","0110001001000XXXXXXXX11","1110001001000XXXXXXXX10","01100010011000111001101","11100010011100111001100","0110001010000XXXXXXXX11","1110001010000XXXXXXXX10","01100010101000111010101","11100010101100111010100","01100010110000111011001","11100010110100111011000","01100010111100111011100","11100010111100111011101","0110001100000XXXXXXXX11","1110001100000XXXXXXXX10","01100011001000111100101","11100011001100111100100","01100011010000111101001","11100011010100111101000","01100011011100111101100","11100011011100111101101","01100011100000111110001","11100011100100111110000","01100011101100111110100","11100011101100111110101","01100011110100111111000","11100011110100111111001","0110001111110XXXXXXXX11","1110001111110XXXXXXXX11","0110010000000XXXXXXXX11","1110010000000XXXXXXXX11","0110010000100XXXXXXXX11","1110010000100XXXXXXXX10","0110010001000XXXXXXXX11","1110010001000XXXXXXXX10","01100100011000110001101","11100100011100110001100","0110010010000XXXXXXXX11","1110010010000XXXXXXXX10","01100100101000110010101","11100100101100110010100","01100100110000110011001","11100100110100110011000","01100100111100110100000","11100100111100110100001","0110010100000XXXXXXXX11","1110010100000XXXXXXXX10","01100101001000110100101","11100101001100110100100","01100101010000110101001","11100101010100110101000","01100101011100110010000","11100101011100110010001","01100101100000110110001","11100101100100110110000","01100101101100110001000","11100101101100110001001","01100101110100110000100","11100101110100110000101","0110010111110XXXXXXXX11","1110010111110XXXXXXXX11","0110011000000XXXXXXXX11","1110011000000XXXXXXXX10","01100110001000111000101","11100110001100111000100","01100110010000111001001","11100110010100111001000","01100110011100111100000","11100110011100111100001","01100110100000111010001","11100110100100111010000","01100110101100111111100","11100110101100111111101","01100110110100111000000","11100110110100111000001","0110011011110XXXXXXXX11","1110011011110XXXXXXXX11","01100111000000110011101","11100111000100110011100","01100111001100110000000","11100111001100110000001","01100111010100110111100","11100111010100110111101","0110011101110XXXXXXXX11","1110011101110XXXXXXXX11","01100111100110111110000","11100111100110111110001","0110011110110XXXXXXXX11","1110011110110XXXXXXXX11","0110011111010XXXXXXXX11","1110011111010XXXXXXXX11","0110011111110XXXXXXXX11","1110011111110XXXXXXXX11","0110100000010XXXXXXXX11","1110100000010XXXXXXXX11","0110100000110XXXXXXXX11","1110100000110XXXXXXXX11","0110100001010XXXXXXXX11","1110100001010XXXXXXXX11","01101000011110001110001","11101000011110001110000","0110100010010XXXXXXXX11","1110100010010XXXXXXXX11","01101000101100000111101","11101000101100000111100","01101000110100000000001","11101000110100000000000","01101000111100000011100","11101000111100000011101","0110100100010XXXXXXXX11","1110100100010XXXXXXXX11","01101001001100001000001","11101001001100001000000","01101001010100001111101","11101001010100001111100","01101001011100000101100","11101001011100000101101","01101001100100001100001","11101001100100001100000","01101001101100000110100","11101001101100000110101","01101001110100000111000","11101001110100000111001","0110100111110XXXXXXXX11","1110100111110XXXXXXXX11","0110101000010XXXXXXXX11","1110101000010XXXXXXXX11","01101010001100000000101","11101010001100000000100","01101010010100000001001","11101010010100000001000","01101010011100001001100","11101010011100001001101","01101010100100000010001","11101010100100000010000","01101010101100001010100","11101010101100001010101","01101010110100001011000","11101010110100001011001","0110101011110XXXXXXXX11","1110101011110XXXXXXXX11","01101011000100000100001","11101011000100000100000","01101011001100001100100","11101011001100001100101","01101011010100001101000","11101011010100001101001","0110101101110XXXXXXXX11","1110101101110XXXXXXXX11","01101011100100001110000","11101011100100001110001","0110101110110XXXXXXXX11","1110101110110XXXXXXXX11","0110101111010XXXXXXXX11","1110101111010XXXXXXXX11","0110101111110XXXXXXXX11","1110101111110XXXXXXXX11","0110110000010XXXXXXXX11","1110110000010XXXXXXXX11","01101100001100001111001","11101100001100001111000","01101100010100001110101","11101100010100001110100","01101100011100000001100","11101100011100000001101","01101100100100001101101","11101100100100001101100","01101100101100000010100","11101100101100000010101","01101100110100000011000","11101100110100000011001","0110110011110XXXXXXXX11","1110110011110XXXXXXXX11","01101101000100001011101","11101101000100001011100","01101101001100000100100","11101101001100000100101","01101101010100000101000","11101101010100000101001","0110110101110XXXXXXXX11","1110110101110XXXXXXXX11","01101101100100000110000","11101101100100000110001","0110110110110XXXXXXXX11","1110110110110XXXXXXXX11","0110110111010XXXXXXXX11","1110110111010XXXXXXXX11","0110110111110XXXXXXXX11","1110110111110XXXXXXXX11","0110111000010XXXXXXXX11","1110111000010XXXXXXXX10","01101110001100001000100","11101110001100001000101","01101110010100001001000","11101110010100001001001","0110111001110XXXXXXXX11","1110111001110XXXXXXXX11","01101110100100001010000","11101110100100001010001","0110111010110XXXXXXXX11","1110111010110XXXXXXXX11","0110111011010XXXXXXXX11","1110111011010XXXXXXXX11","0110111011110XXXXXXXX11","1110111011110XXXXXXXX11","0110111100010XXXXXXXX10","1110111100010XXXXXXXX11","0110111100110XXXXXXXX11","1110111100110XXXXXXXX11","0110111101010XXXXXXXX11","1110111101010XXXXXXXX11","0110111101110XXXXXXXX11","1110111101110XXXXXXXX11","0110111110010XXXXXXXX11","1110111110010XXXXXXXX11","0110111110110XXXXXXXX11","1110111110110XXXXXXXX11","0110111111010XXXXXXXX11","1110111111010XXXXXXXX11","0110111111110XXXXXXXX11","1110111111110XXXXXXXX11","0111000000010XXXXXXXX11","1111000000010XXXXXXXX11","0111000000110XXXXXXXX11","1111000000110XXXXXXXX11","0111000001010XXXXXXXX11","1111000001010XXXXXXXX11","01110000011111111110001","11110000011111111110000","0111000010010XXXXXXXX11","1111000010010XXXXXXXX11","0111000010110XXXXXXXX11","1111000010110XXXXXXXX10","0111000011010XXXXXXXX11","1111000011010XXXXXXXX10","0111000011110XXXXXXXX10","1111000011110XXXXXXXX11","0111000100010XXXXXXXX11","1111000100010XXXXXXXX11","0111000100110XXXXXXXX11","1111000100110XXXXXXXX10","0111000101010XXXXXXXX11","1111000101010XXXXXXXX10","0111000101110XXXXXXXX10","1111000101110XXXXXXXX11","0111000110010XXXXXXXX11","1111000110010XXXXXXXX10","0111000110110XXXXXXXX10","1111000110110XXXXXXXX11","0111000111010XXXXXXXX10","1111000111010XXXXXXXX11","0111000111110XXXXXXXX11","1111000111110XXXXXXXX11","0111001000010XXXXXXXX11","1111001000010XXXXXXXX11","0111001000110XXXXXXXX11","1111001000110XXXXXXXX10","0111001001010XXXXXXXX11","1111001001010XXXXXXXX10","0111001001110XXXXXXXX10","1111001001110XXXXXXXX11","0111001010010XXXXXXXX11","1111001010010XXXXXXXX10","0111001010110XXXXXXXX10","1111001010110XXXXXXXX11","0111001011010XXXXXXXX10","1111001011010XXXXXXXX11","0111001011110XXXXXXXX11","1111001011110XXXXXXXX11","0111001100010XXXXXXXX11","1111001100010XXXXXXXX10","0111001100110XXXXXXXX10","1111001100110XXXXXXXX11","0111001101010XXXXXXXX10","1111001101010XXXXXXXX11","0111001101110XXXXXXXX11","1111001101110XXXXXXXX11","0111001110010XXXXXXXX10","1111001110010XXXXXXXX11","0111001110110XXXXXXXX11","1111001110110XXXXXXXX11","0111001111010XXXXXXXX11","1111001111010XXXXXXXX11","0111001111110XXXXXXXX11","1111001111110XXXXXXXX11","0111010000010XXXXXXXX11","1111010000010XXXXXXXX11","01110100001111111111001","11110100001111111111000","01110100010111111110101","11110100010111111110100","0111010001110XXXXXXXX10","1111010001110XXXXXXXX11","01110100100111111101101","11110100100111111101100","0111010010110XXXXXXXX10","1111010010110XXXXXXXX11","0111010011010XXXXXXXX10","1111010011010XXXXXXXX11","0111010011110XXXXXXXX11","1111010011110XXXXXXXX11","01110101000111111011101","11110101000111111011100","0111010100110XXXXXXXX10","1111010100110XXXXXXXX11","0111010101010XXXXXXXX10","1111010101010XXXXXXXX11","0111010101110XXXXXXXX11","1111010101110XXXXXXXX11","0111010110010XXXXXXXX10","1111010110010XXXXXXXX11","0111010110110XXXXXXXX11","1111010110110XXXXXXXX11","0111010111010XXXXXXXX11","1111010111010XXXXXXXX11","0111010111110XXXXXXXX11","1111010111110XXXXXXXX11","0111011000010XXXXXXXX11","1111011000010XXXXXXXX10","01110110001101111000100","11110110001101111000101","01110110010101111001000","11110110010101111001001","0111011001110XXXXXXXX11","1111011001110XXXXXXXX11","01110110100101111010000","11110110100101111010001","0111011010110XXXXXXXX11","1111011010110XXXXXXXX11","0111011011010XXXXXXXX11","1111011011010XXXXXXXX11","0111011011110XXXXXXXX11","1111011011110XXXXXXXX11","0111011100010XXXXXXXX10","1111011100010XXXXXXXX11","0111011100110XXXXXXXX11","1111011100110XXXXXXXX11","0111011101010XXXXXXXX11","1111011101010XXXXXXXX11","0111011101110XXXXXXXX11","1111011101110XXXXXXXX11","0111011110010XXXXXXXX11","1111011110010XXXXXXXX11","0111011110110XXXXXXXX11","1111011110110XXXXXXXX11","0111011111010XXXXXXXX11","1111011111010XXXXXXXX11","0111011111110XXXXXXXX11","1111011111110XXXXXXXX11","0111100000010XXXXXXXX11","1111100000010XXXXXXXX11","0111100000110XXXXXXXX11","1111100000110XXXXXXXX11","0111100001010XXXXXXXX11","1111100001010XXXXXXXX11","0111100001110XXXXXXXX11","1111100001110XXXXXXXX11","0111100010010XXXXXXXX11","1111100010010XXXXXXXX11","0111100010110XXXXXXXX11","1111100010110XXXXXXXX11","0111100011010XXXXXXXX11","1111100011010XXXXXXXX11","0111100011110XXXXXXXX11","1111100011110XXXXXXXX11","0111100100010XXXXXXXX11","1111100100010XXXXXXXX11","0111100100110XXXXXXXX11","1111100100110XXXXXXXX11","0111100101010XXXXXXXX11","1111100101010XXXXXXXX11","0111100101110XXXXXXXX11","1111100101110XXXXXXXX11","0111100110010XXXXXXXX11","1111100110010XXXXXXXX11","0111100110110XXXXXXXX11","1111100110110XXXXXXXX11","0111100111010XXXXXXXX11","1111100111010XXXXXXXX11","0111100111110XXXXXXXX11","1111100111110XXXXXXXX11","0111101000010XXXXXXXX11","1111101000010XXXXXXXX11","0111101000110XXXXXXXX11","1111101000110XXXXXXXX11","0111101001010XXXXXXXX11","1111101001010XXXXXXXX11","0111101001110XXXXXXXX11","1111101001110XXXXXXXX11","0111101010010XXXXXXXX11","1111101010010XXXXXXXX11","0111101010110XXXXXXXX11","1111101010110XXXXXXXX11","0111101011010XXXXXXXX11","1111101011010XXXXXXXX11","0111101011110XXXXXXXX11","1111101011110XXXXXXXX11","0111101100010XXXXXXXX11","1111101100010XXXXXXXX11","0111101100110XXXXXXXX11","1111101100110XXXXXXXX11","0111101101010XXXXXXXX11","1111101101010XXXXXXXX11","0111101101110XXXXXXXX11","1111101101110XXXXXXXX11","0111101110010XXXXXXXX11","1111101110010XXXXXXXX11","0111101110110XXXXXXXX11","1111101110110XXXXXXXX11","0111101111010XXXXXXXX11","1111101111010XXXXXXXX11","0111101111110XXXXXXXX11","1111101111110XXXXXXXX11","0111110000010XXXXXXXX11","1111110000010XXXXXXXX11","0111110000110XXXXXXXX11","1111110000110XXXXXXXX11","0111110001010XXXXXXXX11","1111110001010XXXXXXXX11","0111110001110XXXXXXXX11","1111110001110XXXXXXXX11","0111110010010XXXXXXXX11","1111110010010XXXXXXXX11","0111110010110XXXXXXXX11","1111110010110XXXXXXXX11","0111110011010XXXXXXXX11","1111110011010XXXXXXXX11","0111110011110XXXXXXXX11","1111110011110XXXXXXXX11","0111110100010XXXXXXXX11","1111110100010XXXXXXXX11","0111110100110XXXXXXXX11","1111110100110XXXXXXXX11","0111110101010XXXXXXXX11","1111110101010XXXXXXXX11","0111110101110XXXXXXXX11","1111110101110XXXXXXXX11","0111110110010XXXXXXXX11","1111110110010XXXXXXXX11","0111110110110XXXXXXXX11","1111110110110XXXXXXXX11","0111110111010XXXXXXXX11","1111110111010XXXXXXXX11","0111110111110XXXXXXXX11","1111110111110XXXXXXXX11","0111111000010XXXXXXXX11","1111111000010XXXXXXXX11","0111111000110XXXXXXXX11","1111111000110XXXXXXXX11","0111111001010XXXXXXXX11","1111111001010XXXXXXXX11","0111111001110XXXXXXXX11","1111111001110XXXXXXXX11","0111111010010XXXXXXXX11","1111111010010XXXXXXXX11","0111111010110XXXXXXXX11","1111111010110XXXXXXXX11","0111111011010XXXXXXXX11","1111111011010XXXXXXXX11","0111111011110XXXXXXXX11","1111111011110XXXXXXXX11","0111111100010XXXXXXXX11","1111111100010XXXXXXXX11","0111111100110XXXXXXXX11","1111111100110XXXXXXXX11","0111111101010XXXXXXXX11","1111111101010XXXXXXXX11","0111111101110XXXXXXXX11","1111111101110XXXXXXXX11","0111111110010XXXXXXXX11","1111111110010XXXXXXXX11","0111111110110XXXXXXXX11","1111111110110XXXXXXXX11","0111111111010XXXXXXXX11","1111111111010XXXXXXXX11","0111111111110XXXXXXXX11","1111111111110XXXXXXXX11",
        others => (others => 'X')
    );

    constant CLK_MHZ : positive := 100;
    signal clk, reset_n : std_logic := '0';

    signal e8b : std_logic_vector(8 downto 0);
    signal e10b : std_logic_vector(9 downto 0);
    signal edin, edout, eerr : std_logic;
    signal d8b : std_logic_vector(8 downto 0);
    signal d10b : std_logic_vector(9 downto 0);
    signal ddin, ddout, dderr, derr : std_logic;

begin

    clk <= not clk after (500 ns / CLK_MHZ);
    reset_n <= '0', '1' after 100 ns;

    i_enc : entity work.enc_8b10b
    port map (
        datain => e8b,
        dispin => edin,
        dataout => e10b,
        dispout => edout,
        err => eerr--,
    );

    i_dec : entity work.dec_8b10b
    port map (
        datain => d10b,
        dispin => ddin,
        dataout => d8b,
        dispout => ddout,
        disperr => dderr,
        err => derr--,
    );

    process
    begin
        wait until rising_edge(reset_n);

        for i in data_enc'range loop
            edin <= data_enc(i)(0);
            e8b <= data_enc(i)(1 to 9);
            wait until rising_edge(clk);
            if ( edout & e10b & eerr /= data_enc(i)(10 to 21) ) then
                report integer'image(i);
                report "edout & e10b & eerr /= " & work.util.to_string(data_enc(i)(10 to 21));
            end if;
        end loop;



        for i in data_dec'range loop
            ddin <= data_dec(i)(0);
            d10b <= data_dec(i)(1 to 10);
            wait until rising_edge(clk);

            assert ( ddout = data_dec(i)(11) ) report "" severity failure;
            assert ( (derr or dderr) = (data_dec(i)(21) or data_dec(i)(22)) ) report "" severity failure;

            if ( derr = '0' and dderr = '0' and data_dec(i)(21 to 22) = "00" ) then
                assert ( ddout & d8b & derr & dderr = data_dec(i)(11 to 22) ) report "" severity failure;
            end if;

            if ( derr = '1' and data_dec(i)(21) = '1' ) then
                --
            elsif ( ddout & d8b & derr & dderr /= data_dec(i)(11 to 22) ) then
                report integer'image(i);
                report work.util.to_string(data_dec(i)(0 to 10)) & " =>                " & work.util.to_string(ddout & d8b & derr & dderr);
                report "ddout & d8b & derr & dderr /= " & work.util.to_string(data_dec(i)(11 to 22));
                report "                              " & work.util.to_string(ddout & d8b & derr & dderr xor data_dec(i)(11 to 22));
            end if;

        end loop;

        wait;
    end process;

end architecture;
